library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

package table_h_package is 
  type table_h is array (0 to 65535) of std_logic_vector(7 downto 0);
constant table : table_h := (  
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 

  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 

  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 

  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 
  x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00",   x"00", 

  x"00",   x"01",   x"02",   x"03",   x"04",   x"05",   x"06",   x"07", 
  x"08",   x"09",   x"0A",   x"0B",   x"0C",   x"0D",   x"0E",   x"0F", 
  x"10",   x"11",   x"12",   x"13",   x"14",   x"15",   x"16",   x"17", 
  x"18",   x"19",   x"1A",   x"1B",   x"1C",   x"1D",   x"1E",   x"1F", 
  x"20",   x"21",   x"22",   x"23",   x"24",   x"25",   x"26",   x"27", 
  x"28",   x"29",   x"2A",   x"2B",   x"2C",   x"2D",   x"2E",   x"2F", 
  x"30",   x"31",   x"32",   x"33",   x"34",   x"35",   x"36",   x"37", 
  x"38",   x"39",   x"3A",   x"3B",   x"3C",   x"3D",   x"3E",   x"3F", 
  x"40",   x"41",   x"42",   x"43",   x"44",   x"45",   x"46",   x"47", 
  x"48",   x"49",   x"4A",   x"4B",   x"4C",   x"4D",   x"4E",   x"4F", 
  x"50",   x"51",   x"52",   x"53",   x"54",   x"55",   x"56",   x"57", 
  x"58",   x"59",   x"5A",   x"5B",   x"5C",   x"5D",   x"5E",   x"5F", 
  x"60",   x"61",   x"62",   x"63",   x"64",   x"65",   x"66",   x"67", 
  x"68",   x"69",   x"6A",   x"6B",   x"6C",   x"6D",   x"6E",   x"6F", 
  x"70",   x"71",   x"72",   x"73",   x"74",   x"75",   x"76",   x"77", 
  x"78",   x"79",   x"7A",   x"7B",   x"7C",   x"7D",   x"7E",   x"7F", 
  x"80",   x"81",   x"82",   x"83",   x"84",   x"85",   x"86",   x"87", 
  x"88",   x"89",   x"8A",   x"8B",   x"8C",   x"8D",   x"8E",   x"8F", 
  x"90",   x"91",   x"92",   x"93",   x"94",   x"95",   x"96",   x"97", 
  x"98",   x"99",   x"9A",   x"9B",   x"9C",   x"9D",   x"9E",   x"9F", 
  x"A0",   x"A1",   x"A2",   x"A3",   x"A4",   x"A5",   x"A6",   x"A7", 
  x"A8",   x"A9",   x"AA",   x"AB",   x"AC",   x"AD",   x"AE",   x"AF", 
  x"B0",   x"B1",   x"B2",   x"B3",   x"B4",   x"B5",   x"B6",   x"B7", 
  x"B8",   x"B9",   x"BA",   x"BB",   x"BC",   x"BD",   x"BE",   x"BF", 
  x"C0",   x"C1",   x"C2",   x"C3",   x"C4",   x"C5",   x"C6",   x"C7", 
  x"C8",   x"C9",   x"CA",   x"CB",   x"CC",   x"CD",   x"CE",   x"CF", 
  x"D0",   x"D1",   x"D2",   x"D3",   x"D4",   x"D5",   x"D6",   x"D7", 
  x"D8",   x"D9",   x"DA",   x"DB",   x"DC",   x"DD",   x"DE",   x"DF", 
  x"E0",   x"E1",   x"E2",   x"E3",   x"E4",   x"E5",   x"E6",   x"E7", 
  x"E8",   x"E9",   x"EA",   x"EB",   x"EC",   x"ED",   x"EE",   x"EF", 
  x"F0",   x"F1",   x"F2",   x"F3",   x"F4",   x"F5",   x"F6",   x"F7", 
  x"F8",   x"F9",   x"FA",   x"FB",   x"FC",   x"FD",   x"FE",   x"FF", 
  x"00",   x"02",   x"04",   x"06",   x"08",   x"0A",   x"0C",   x"0E", 
  x"10",   x"12",   x"14",   x"16",   x"18",   x"1A",   x"1C",   x"1E", 
  x"20",   x"22",   x"24",   x"26",   x"28",   x"2A",   x"2C",   x"2E", 
  x"30",   x"32",   x"34",   x"36",   x"38",   x"3A",   x"3C",   x"3E", 
  x"40",   x"42",   x"44",   x"46",   x"48",   x"4A",   x"4C",   x"4E", 
  x"50",   x"52",   x"54",   x"56",   x"58",   x"5A",   x"5C",   x"5E", 
  x"60",   x"62",   x"64",   x"66",   x"68",   x"6A",   x"6C",   x"6E", 
  x"70",   x"72",   x"74",   x"76",   x"78",   x"7A",   x"7C",   x"7E", 
  x"80",   x"82",   x"84",   x"86",   x"88",   x"8A",   x"8C",   x"8E", 
  x"90",   x"92",   x"94",   x"96",   x"98",   x"9A",   x"9C",   x"9E", 
  x"A0",   x"A2",   x"A4",   x"A6",   x"A8",   x"AA",   x"AC",   x"AE", 
  x"B0",   x"B2",   x"B4",   x"B6",   x"B8",   x"BA",   x"BC",   x"BE", 
  x"C0",   x"C2",   x"C4",   x"C6",   x"C8",   x"CA",   x"CC",   x"CE", 
  x"D0",   x"D2",   x"D4",   x"D6",   x"D8",   x"DA",   x"DC",   x"DE", 
  x"E0",   x"E2",   x"E4",   x"E6",   x"E8",   x"EA",   x"EC",   x"EE", 
  x"F0",   x"F2",   x"F4",   x"F6",   x"F8",   x"FA",   x"FC",   x"FE", 
  x"C3",   x"C1",   x"C7",   x"C5",   x"CB",   x"C9",   x"CF",   x"CD", 
  x"D3",   x"D1",   x"D7",   x"D5",   x"DB",   x"D9",   x"DF",   x"DD", 
  x"E3",   x"E1",   x"E7",   x"E5",   x"EB",   x"E9",   x"EF",   x"ED", 
  x"F3",   x"F1",   x"F7",   x"F5",   x"FB",   x"F9",   x"FF",   x"FD", 
  x"83",   x"81",   x"87",   x"85",   x"8B",   x"89",   x"8F",   x"8D", 
  x"93",   x"91",   x"97",   x"95",   x"9B",   x"99",   x"9F",   x"9D", 
  x"A3",   x"A1",   x"A7",   x"A5",   x"AB",   x"A9",   x"AF",   x"AD", 
  x"B3",   x"B1",   x"B7",   x"B5",   x"BB",   x"B9",   x"BF",   x"BD", 
  x"43",   x"41",   x"47",   x"45",   x"4B",   x"49",   x"4F",   x"4D", 
  x"53",   x"51",   x"57",   x"55",   x"5B",   x"59",   x"5F",   x"5D", 
  x"63",   x"61",   x"67",   x"65",   x"6B",   x"69",   x"6F",   x"6D", 
  x"73",   x"71",   x"77",   x"75",   x"7B",   x"79",   x"7F",   x"7D", 
  x"03",   x"01",   x"07",   x"05",   x"0B",   x"09",   x"0F",   x"0D", 
  x"13",   x"11",   x"17",   x"15",   x"1B",   x"19",   x"1F",   x"1D", 
  x"23",   x"21",   x"27",   x"25",   x"2B",   x"29",   x"2F",   x"2D", 
  x"33",   x"31",   x"37",   x"35",   x"3B",   x"39",   x"3F",   x"3D", 
  x"00",   x"03",   x"06",   x"05",   x"0C",   x"0F",   x"0A",   x"09", 
  x"18",   x"1B",   x"1E",   x"1D",   x"14",   x"17",   x"12",   x"11", 
  x"30",   x"33",   x"36",   x"35",   x"3C",   x"3F",   x"3A",   x"39", 
  x"28",   x"2B",   x"2E",   x"2D",   x"24",   x"27",   x"22",   x"21", 
  x"60",   x"63",   x"66",   x"65",   x"6C",   x"6F",   x"6A",   x"69", 
  x"78",   x"7B",   x"7E",   x"7D",   x"74",   x"77",   x"72",   x"71", 
  x"50",   x"53",   x"56",   x"55",   x"5C",   x"5F",   x"5A",   x"59", 
  x"48",   x"4B",   x"4E",   x"4D",   x"44",   x"47",   x"42",   x"41", 
  x"C0",   x"C3",   x"C6",   x"C5",   x"CC",   x"CF",   x"CA",   x"C9", 
  x"D8",   x"DB",   x"DE",   x"DD",   x"D4",   x"D7",   x"D2",   x"D1", 
  x"F0",   x"F3",   x"F6",   x"F5",   x"FC",   x"FF",   x"FA",   x"F9", 
  x"E8",   x"EB",   x"EE",   x"ED",   x"E4",   x"E7",   x"E2",   x"E1", 
  x"A0",   x"A3",   x"A6",   x"A5",   x"AC",   x"AF",   x"AA",   x"A9", 
  x"B8",   x"BB",   x"BE",   x"BD",   x"B4",   x"B7",   x"B2",   x"B1", 
  x"90",   x"93",   x"96",   x"95",   x"9C",   x"9F",   x"9A",   x"99", 
  x"88",   x"8B",   x"8E",   x"8D",   x"84",   x"87",   x"82",   x"81", 
  x"43",   x"40",   x"45",   x"46",   x"4F",   x"4C",   x"49",   x"4A", 
  x"5B",   x"58",   x"5D",   x"5E",   x"57",   x"54",   x"51",   x"52", 
  x"73",   x"70",   x"75",   x"76",   x"7F",   x"7C",   x"79",   x"7A", 
  x"6B",   x"68",   x"6D",   x"6E",   x"67",   x"64",   x"61",   x"62", 
  x"23",   x"20",   x"25",   x"26",   x"2F",   x"2C",   x"29",   x"2A", 
  x"3B",   x"38",   x"3D",   x"3E",   x"37",   x"34",   x"31",   x"32", 
  x"13",   x"10",   x"15",   x"16",   x"1F",   x"1C",   x"19",   x"1A", 
  x"0B",   x"08",   x"0D",   x"0E",   x"07",   x"04",   x"01",   x"02", 
  x"83",   x"80",   x"85",   x"86",   x"8F",   x"8C",   x"89",   x"8A", 
  x"9B",   x"98",   x"9D",   x"9E",   x"97",   x"94",   x"91",   x"92", 
  x"B3",   x"B0",   x"B5",   x"B6",   x"BF",   x"BC",   x"B9",   x"BA", 
  x"AB",   x"A8",   x"AD",   x"AE",   x"A7",   x"A4",   x"A1",   x"A2", 
  x"E3",   x"E0",   x"E5",   x"E6",   x"EF",   x"EC",   x"E9",   x"EA", 
  x"FB",   x"F8",   x"FD",   x"FE",   x"F7",   x"F4",   x"F1",   x"F2", 
  x"D3",   x"D0",   x"D5",   x"D6",   x"DF",   x"DC",   x"D9",   x"DA", 
  x"CB",   x"C8",   x"CD",   x"CE",   x"C7",   x"C4",   x"C1",   x"C2", 
  x"00",   x"04",   x"08",   x"0C",   x"10",   x"14",   x"18",   x"1C", 
  x"20",   x"24",   x"28",   x"2C",   x"30",   x"34",   x"38",   x"3C", 
  x"40",   x"44",   x"48",   x"4C",   x"50",   x"54",   x"58",   x"5C", 
  x"60",   x"64",   x"68",   x"6C",   x"70",   x"74",   x"78",   x"7C", 
  x"80",   x"84",   x"88",   x"8C",   x"90",   x"94",   x"98",   x"9C", 
  x"A0",   x"A4",   x"A8",   x"AC",   x"B0",   x"B4",   x"B8",   x"BC", 
  x"C0",   x"C4",   x"C8",   x"CC",   x"D0",   x"D4",   x"D8",   x"DC", 
  x"E0",   x"E4",   x"E8",   x"EC",   x"F0",   x"F4",   x"F8",   x"FC", 
  x"C3",   x"C7",   x"CB",   x"CF",   x"D3",   x"D7",   x"DB",   x"DF", 
  x"E3",   x"E7",   x"EB",   x"EF",   x"F3",   x"F7",   x"FB",   x"FF", 
  x"83",   x"87",   x"8B",   x"8F",   x"93",   x"97",   x"9B",   x"9F", 
  x"A3",   x"A7",   x"AB",   x"AF",   x"B3",   x"B7",   x"BB",   x"BF", 
  x"43",   x"47",   x"4B",   x"4F",   x"53",   x"57",   x"5B",   x"5F", 
  x"63",   x"67",   x"6B",   x"6F",   x"73",   x"77",   x"7B",   x"7F", 
  x"03",   x"07",   x"0B",   x"0F",   x"13",   x"17",   x"1B",   x"1F", 
  x"23",   x"27",   x"2B",   x"2F",   x"33",   x"37",   x"3B",   x"3F", 
  x"45",   x"41",   x"4D",   x"49",   x"55",   x"51",   x"5D",   x"59", 
  x"65",   x"61",   x"6D",   x"69",   x"75",   x"71",   x"7D",   x"79", 
  x"05",   x"01",   x"0D",   x"09",   x"15",   x"11",   x"1D",   x"19", 
  x"25",   x"21",   x"2D",   x"29",   x"35",   x"31",   x"3D",   x"39", 
  x"C5",   x"C1",   x"CD",   x"C9",   x"D5",   x"D1",   x"DD",   x"D9", 
  x"E5",   x"E1",   x"ED",   x"E9",   x"F5",   x"F1",   x"FD",   x"F9", 
  x"85",   x"81",   x"8D",   x"89",   x"95",   x"91",   x"9D",   x"99", 
  x"A5",   x"A1",   x"AD",   x"A9",   x"B5",   x"B1",   x"BD",   x"B9", 
  x"86",   x"82",   x"8E",   x"8A",   x"96",   x"92",   x"9E",   x"9A", 
  x"A6",   x"A2",   x"AE",   x"AA",   x"B6",   x"B2",   x"BE",   x"BA", 
  x"C6",   x"C2",   x"CE",   x"CA",   x"D6",   x"D2",   x"DE",   x"DA", 
  x"E6",   x"E2",   x"EE",   x"EA",   x"F6",   x"F2",   x"FE",   x"FA", 
  x"06",   x"02",   x"0E",   x"0A",   x"16",   x"12",   x"1E",   x"1A", 
  x"26",   x"22",   x"2E",   x"2A",   x"36",   x"32",   x"3E",   x"3A", 
  x"46",   x"42",   x"4E",   x"4A",   x"56",   x"52",   x"5E",   x"5A", 
  x"66",   x"62",   x"6E",   x"6A",   x"76",   x"72",   x"7E",   x"7A", 
  x"00",   x"05",   x"0A",   x"0F",   x"14",   x"11",   x"1E",   x"1B", 
  x"28",   x"2D",   x"22",   x"27",   x"3C",   x"39",   x"36",   x"33", 
  x"50",   x"55",   x"5A",   x"5F",   x"44",   x"41",   x"4E",   x"4B", 
  x"78",   x"7D",   x"72",   x"77",   x"6C",   x"69",   x"66",   x"63", 
  x"A0",   x"A5",   x"AA",   x"AF",   x"B4",   x"B1",   x"BE",   x"BB", 
  x"88",   x"8D",   x"82",   x"87",   x"9C",   x"99",   x"96",   x"93", 
  x"F0",   x"F5",   x"FA",   x"FF",   x"E4",   x"E1",   x"EE",   x"EB", 
  x"D8",   x"DD",   x"D2",   x"D7",   x"CC",   x"C9",   x"C6",   x"C3", 
  x"83",   x"86",   x"89",   x"8C",   x"97",   x"92",   x"9D",   x"98", 
  x"AB",   x"AE",   x"A1",   x"A4",   x"BF",   x"BA",   x"B5",   x"B0", 
  x"D3",   x"D6",   x"D9",   x"DC",   x"C7",   x"C2",   x"CD",   x"C8", 
  x"FB",   x"FE",   x"F1",   x"F4",   x"EF",   x"EA",   x"E5",   x"E0", 
  x"23",   x"26",   x"29",   x"2C",   x"37",   x"32",   x"3D",   x"38", 
  x"0B",   x"0E",   x"01",   x"04",   x"1F",   x"1A",   x"15",   x"10", 
  x"73",   x"76",   x"79",   x"7C",   x"67",   x"62",   x"6D",   x"68", 
  x"5B",   x"5E",   x"51",   x"54",   x"4F",   x"4A",   x"45",   x"40", 
  x"C5",   x"C0",   x"CF",   x"CA",   x"D1",   x"D4",   x"DB",   x"DE", 
  x"ED",   x"E8",   x"E7",   x"E2",   x"F9",   x"FC",   x"F3",   x"F6", 
  x"95",   x"90",   x"9F",   x"9A",   x"81",   x"84",   x"8B",   x"8E", 
  x"BD",   x"B8",   x"B7",   x"B2",   x"A9",   x"AC",   x"A3",   x"A6", 
  x"65",   x"60",   x"6F",   x"6A",   x"71",   x"74",   x"7B",   x"7E", 
  x"4D",   x"48",   x"47",   x"42",   x"59",   x"5C",   x"53",   x"56", 
  x"35",   x"30",   x"3F",   x"3A",   x"21",   x"24",   x"2B",   x"2E", 
  x"1D",   x"18",   x"17",   x"12",   x"09",   x"0C",   x"03",   x"06", 
  x"46",   x"43",   x"4C",   x"49",   x"52",   x"57",   x"58",   x"5D", 
  x"6E",   x"6B",   x"64",   x"61",   x"7A",   x"7F",   x"70",   x"75", 
  x"16",   x"13",   x"1C",   x"19",   x"02",   x"07",   x"08",   x"0D", 
  x"3E",   x"3B",   x"34",   x"31",   x"2A",   x"2F",   x"20",   x"25", 
  x"E6",   x"E3",   x"EC",   x"E9",   x"F2",   x"F7",   x"F8",   x"FD", 
  x"CE",   x"CB",   x"C4",   x"C1",   x"DA",   x"DF",   x"D0",   x"D5", 
  x"B6",   x"B3",   x"BC",   x"B9",   x"A2",   x"A7",   x"A8",   x"AD", 
  x"9E",   x"9B",   x"94",   x"91",   x"8A",   x"8F",   x"80",   x"85", 
  x"00",   x"06",   x"0C",   x"0A",   x"18",   x"1E",   x"14",   x"12", 
  x"30",   x"36",   x"3C",   x"3A",   x"28",   x"2E",   x"24",   x"22", 
  x"60",   x"66",   x"6C",   x"6A",   x"78",   x"7E",   x"74",   x"72", 
  x"50",   x"56",   x"5C",   x"5A",   x"48",   x"4E",   x"44",   x"42", 
  x"C0",   x"C6",   x"CC",   x"CA",   x"D8",   x"DE",   x"D4",   x"D2", 
  x"F0",   x"F6",   x"FC",   x"FA",   x"E8",   x"EE",   x"E4",   x"E2", 
  x"A0",   x"A6",   x"AC",   x"AA",   x"B8",   x"BE",   x"B4",   x"B2", 
  x"90",   x"96",   x"9C",   x"9A",   x"88",   x"8E",   x"84",   x"82", 
  x"43",   x"45",   x"4F",   x"49",   x"5B",   x"5D",   x"57",   x"51", 
  x"73",   x"75",   x"7F",   x"79",   x"6B",   x"6D",   x"67",   x"61", 
  x"23",   x"25",   x"2F",   x"29",   x"3B",   x"3D",   x"37",   x"31", 
  x"13",   x"15",   x"1F",   x"19",   x"0B",   x"0D",   x"07",   x"01", 
  x"83",   x"85",   x"8F",   x"89",   x"9B",   x"9D",   x"97",   x"91", 
  x"B3",   x"B5",   x"BF",   x"B9",   x"AB",   x"AD",   x"A7",   x"A1", 
  x"E3",   x"E5",   x"EF",   x"E9",   x"FB",   x"FD",   x"F7",   x"F1", 
  x"D3",   x"D5",   x"DF",   x"D9",   x"CB",   x"CD",   x"C7",   x"C1", 
  x"86",   x"80",   x"8A",   x"8C",   x"9E",   x"98",   x"92",   x"94", 
  x"B6",   x"B0",   x"BA",   x"BC",   x"AE",   x"A8",   x"A2",   x"A4", 
  x"E6",   x"E0",   x"EA",   x"EC",   x"FE",   x"F8",   x"F2",   x"F4", 
  x"D6",   x"D0",   x"DA",   x"DC",   x"CE",   x"C8",   x"C2",   x"C4", 
  x"46",   x"40",   x"4A",   x"4C",   x"5E",   x"58",   x"52",   x"54", 
  x"76",   x"70",   x"7A",   x"7C",   x"6E",   x"68",   x"62",   x"64", 
  x"26",   x"20",   x"2A",   x"2C",   x"3E",   x"38",   x"32",   x"34", 
  x"16",   x"10",   x"1A",   x"1C",   x"0E",   x"08",   x"02",   x"04", 
  x"C5",   x"C3",   x"C9",   x"CF",   x"DD",   x"DB",   x"D1",   x"D7", 
  x"F5",   x"F3",   x"F9",   x"FF",   x"ED",   x"EB",   x"E1",   x"E7", 
  x"A5",   x"A3",   x"A9",   x"AF",   x"BD",   x"BB",   x"B1",   x"B7", 
  x"95",   x"93",   x"99",   x"9F",   x"8D",   x"8B",   x"81",   x"87", 
  x"05",   x"03",   x"09",   x"0F",   x"1D",   x"1B",   x"11",   x"17", 
  x"35",   x"33",   x"39",   x"3F",   x"2D",   x"2B",   x"21",   x"27", 
  x"65",   x"63",   x"69",   x"6F",   x"7D",   x"7B",   x"71",   x"77", 
  x"55",   x"53",   x"59",   x"5F",   x"4D",   x"4B",   x"41",   x"47", 
  x"00",   x"07",   x"0E",   x"09",   x"1C",   x"1B",   x"12",   x"15", 
  x"38",   x"3F",   x"36",   x"31",   x"24",   x"23",   x"2A",   x"2D", 
  x"70",   x"77",   x"7E",   x"79",   x"6C",   x"6B",   x"62",   x"65", 
  x"48",   x"4F",   x"46",   x"41",   x"54",   x"53",   x"5A",   x"5D", 
  x"E0",   x"E7",   x"EE",   x"E9",   x"FC",   x"FB",   x"F2",   x"F5", 
  x"D8",   x"DF",   x"D6",   x"D1",   x"C4",   x"C3",   x"CA",   x"CD", 
  x"90",   x"97",   x"9E",   x"99",   x"8C",   x"8B",   x"82",   x"85", 
  x"A8",   x"AF",   x"A6",   x"A1",   x"B4",   x"B3",   x"BA",   x"BD", 
  x"03",   x"04",   x"0D",   x"0A",   x"1F",   x"18",   x"11",   x"16", 
  x"3B",   x"3C",   x"35",   x"32",   x"27",   x"20",   x"29",   x"2E", 
  x"73",   x"74",   x"7D",   x"7A",   x"6F",   x"68",   x"61",   x"66", 
  x"4B",   x"4C",   x"45",   x"42",   x"57",   x"50",   x"59",   x"5E", 
  x"E3",   x"E4",   x"ED",   x"EA",   x"FF",   x"F8",   x"F1",   x"F6", 
  x"DB",   x"DC",   x"D5",   x"D2",   x"C7",   x"C0",   x"C9",   x"CE", 
  x"93",   x"94",   x"9D",   x"9A",   x"8F",   x"88",   x"81",   x"86", 
  x"AB",   x"AC",   x"A5",   x"A2",   x"B7",   x"B0",   x"B9",   x"BE", 
  x"06",   x"01",   x"08",   x"0F",   x"1A",   x"1D",   x"14",   x"13", 
  x"3E",   x"39",   x"30",   x"37",   x"22",   x"25",   x"2C",   x"2B", 
  x"76",   x"71",   x"78",   x"7F",   x"6A",   x"6D",   x"64",   x"63", 
  x"4E",   x"49",   x"40",   x"47",   x"52",   x"55",   x"5C",   x"5B", 
  x"E6",   x"E1",   x"E8",   x"EF",   x"FA",   x"FD",   x"F4",   x"F3", 
  x"DE",   x"D9",   x"D0",   x"D7",   x"C2",   x"C5",   x"CC",   x"CB", 
  x"96",   x"91",   x"98",   x"9F",   x"8A",   x"8D",   x"84",   x"83", 
  x"AE",   x"A9",   x"A0",   x"A7",   x"B2",   x"B5",   x"BC",   x"BB", 
  x"05",   x"02",   x"0B",   x"0C",   x"19",   x"1E",   x"17",   x"10", 
  x"3D",   x"3A",   x"33",   x"34",   x"21",   x"26",   x"2F",   x"28", 
  x"75",   x"72",   x"7B",   x"7C",   x"69",   x"6E",   x"67",   x"60", 
  x"4D",   x"4A",   x"43",   x"44",   x"51",   x"56",   x"5F",   x"58", 
  x"E5",   x"E2",   x"EB",   x"EC",   x"F9",   x"FE",   x"F7",   x"F0", 
  x"DD",   x"DA",   x"D3",   x"D4",   x"C1",   x"C6",   x"CF",   x"C8", 
  x"95",   x"92",   x"9B",   x"9C",   x"89",   x"8E",   x"87",   x"80", 
  x"AD",   x"AA",   x"A3",   x"A4",   x"B1",   x"B6",   x"BF",   x"B8", 
  x"00",   x"08",   x"10",   x"18",   x"20",   x"28",   x"30",   x"38", 
  x"40",   x"48",   x"50",   x"58",   x"60",   x"68",   x"70",   x"78", 
  x"80",   x"88",   x"90",   x"98",   x"A0",   x"A8",   x"B0",   x"B8", 
  x"C0",   x"C8",   x"D0",   x"D8",   x"E0",   x"E8",   x"F0",   x"F8", 
  x"C3",   x"CB",   x"D3",   x"DB",   x"E3",   x"EB",   x"F3",   x"FB", 
  x"83",   x"8B",   x"93",   x"9B",   x"A3",   x"AB",   x"B3",   x"BB", 
  x"43",   x"4B",   x"53",   x"5B",   x"63",   x"6B",   x"73",   x"7B", 
  x"03",   x"0B",   x"13",   x"1B",   x"23",   x"2B",   x"33",   x"3B", 
  x"45",   x"4D",   x"55",   x"5D",   x"65",   x"6D",   x"75",   x"7D", 
  x"05",   x"0D",   x"15",   x"1D",   x"25",   x"2D",   x"35",   x"3D", 
  x"C5",   x"CD",   x"D5",   x"DD",   x"E5",   x"ED",   x"F5",   x"FD", 
  x"85",   x"8D",   x"95",   x"9D",   x"A5",   x"AD",   x"B5",   x"BD", 
  x"86",   x"8E",   x"96",   x"9E",   x"A6",   x"AE",   x"B6",   x"BE", 
  x"C6",   x"CE",   x"D6",   x"DE",   x"E6",   x"EE",   x"F6",   x"FE", 
  x"06",   x"0E",   x"16",   x"1E",   x"26",   x"2E",   x"36",   x"3E", 
  x"46",   x"4E",   x"56",   x"5E",   x"66",   x"6E",   x"76",   x"7E", 
  x"8A",   x"82",   x"9A",   x"92",   x"AA",   x"A2",   x"BA",   x"B2", 
  x"CA",   x"C2",   x"DA",   x"D2",   x"EA",   x"E2",   x"FA",   x"F2", 
  x"0A",   x"02",   x"1A",   x"12",   x"2A",   x"22",   x"3A",   x"32", 
  x"4A",   x"42",   x"5A",   x"52",   x"6A",   x"62",   x"7A",   x"72", 
  x"49",   x"41",   x"59",   x"51",   x"69",   x"61",   x"79",   x"71", 
  x"09",   x"01",   x"19",   x"11",   x"29",   x"21",   x"39",   x"31", 
  x"C9",   x"C1",   x"D9",   x"D1",   x"E9",   x"E1",   x"F9",   x"F1", 
  x"89",   x"81",   x"99",   x"91",   x"A9",   x"A1",   x"B9",   x"B1", 
  x"CF",   x"C7",   x"DF",   x"D7",   x"EF",   x"E7",   x"FF",   x"F7", 
  x"8F",   x"87",   x"9F",   x"97",   x"AF",   x"A7",   x"BF",   x"B7", 
  x"4F",   x"47",   x"5F",   x"57",   x"6F",   x"67",   x"7F",   x"77", 
  x"0F",   x"07",   x"1F",   x"17",   x"2F",   x"27",   x"3F",   x"37", 
  x"0C",   x"04",   x"1C",   x"14",   x"2C",   x"24",   x"3C",   x"34", 
  x"4C",   x"44",   x"5C",   x"54",   x"6C",   x"64",   x"7C",   x"74", 
  x"8C",   x"84",   x"9C",   x"94",   x"AC",   x"A4",   x"BC",   x"B4", 
  x"CC",   x"C4",   x"DC",   x"D4",   x"EC",   x"E4",   x"FC",   x"F4", 
  x"00",   x"09",   x"12",   x"1B",   x"24",   x"2D",   x"36",   x"3F", 
  x"48",   x"41",   x"5A",   x"53",   x"6C",   x"65",   x"7E",   x"77", 
  x"90",   x"99",   x"82",   x"8B",   x"B4",   x"BD",   x"A6",   x"AF", 
  x"D8",   x"D1",   x"CA",   x"C3",   x"FC",   x"F5",   x"EE",   x"E7", 
  x"E3",   x"EA",   x"F1",   x"F8",   x"C7",   x"CE",   x"D5",   x"DC", 
  x"AB",   x"A2",   x"B9",   x"B0",   x"8F",   x"86",   x"9D",   x"94", 
  x"73",   x"7A",   x"61",   x"68",   x"57",   x"5E",   x"45",   x"4C", 
  x"3B",   x"32",   x"29",   x"20",   x"1F",   x"16",   x"0D",   x"04", 
  x"05",   x"0C",   x"17",   x"1E",   x"21",   x"28",   x"33",   x"3A", 
  x"4D",   x"44",   x"5F",   x"56",   x"69",   x"60",   x"7B",   x"72", 
  x"95",   x"9C",   x"87",   x"8E",   x"B1",   x"B8",   x"A3",   x"AA", 
  x"DD",   x"D4",   x"CF",   x"C6",   x"F9",   x"F0",   x"EB",   x"E2", 
  x"E6",   x"EF",   x"F4",   x"FD",   x"C2",   x"CB",   x"D0",   x"D9", 
  x"AE",   x"A7",   x"BC",   x"B5",   x"8A",   x"83",   x"98",   x"91", 
  x"76",   x"7F",   x"64",   x"6D",   x"52",   x"5B",   x"40",   x"49", 
  x"3E",   x"37",   x"2C",   x"25",   x"1A",   x"13",   x"08",   x"01", 
  x"0A",   x"03",   x"18",   x"11",   x"2E",   x"27",   x"3C",   x"35", 
  x"42",   x"4B",   x"50",   x"59",   x"66",   x"6F",   x"74",   x"7D", 
  x"9A",   x"93",   x"88",   x"81",   x"BE",   x"B7",   x"AC",   x"A5", 
  x"D2",   x"DB",   x"C0",   x"C9",   x"F6",   x"FF",   x"E4",   x"ED", 
  x"E9",   x"E0",   x"FB",   x"F2",   x"CD",   x"C4",   x"DF",   x"D6", 
  x"A1",   x"A8",   x"B3",   x"BA",   x"85",   x"8C",   x"97",   x"9E", 
  x"79",   x"70",   x"6B",   x"62",   x"5D",   x"54",   x"4F",   x"46", 
  x"31",   x"38",   x"23",   x"2A",   x"15",   x"1C",   x"07",   x"0E", 
  x"0F",   x"06",   x"1D",   x"14",   x"2B",   x"22",   x"39",   x"30", 
  x"47",   x"4E",   x"55",   x"5C",   x"63",   x"6A",   x"71",   x"78", 
  x"9F",   x"96",   x"8D",   x"84",   x"BB",   x"B2",   x"A9",   x"A0", 
  x"D7",   x"DE",   x"C5",   x"CC",   x"F3",   x"FA",   x"E1",   x"E8", 
  x"EC",   x"E5",   x"FE",   x"F7",   x"C8",   x"C1",   x"DA",   x"D3", 
  x"A4",   x"AD",   x"B6",   x"BF",   x"80",   x"89",   x"92",   x"9B", 
  x"7C",   x"75",   x"6E",   x"67",   x"58",   x"51",   x"4A",   x"43", 
  x"34",   x"3D",   x"26",   x"2F",   x"10",   x"19",   x"02",   x"0B", 
  x"00",   x"0A",   x"14",   x"1E",   x"28",   x"22",   x"3C",   x"36", 
  x"50",   x"5A",   x"44",   x"4E",   x"78",   x"72",   x"6C",   x"66", 
  x"A0",   x"AA",   x"B4",   x"BE",   x"88",   x"82",   x"9C",   x"96", 
  x"F0",   x"FA",   x"E4",   x"EE",   x"D8",   x"D2",   x"CC",   x"C6", 
  x"83",   x"89",   x"97",   x"9D",   x"AB",   x"A1",   x"BF",   x"B5", 
  x"D3",   x"D9",   x"C7",   x"CD",   x"FB",   x"F1",   x"EF",   x"E5", 
  x"23",   x"29",   x"37",   x"3D",   x"0B",   x"01",   x"1F",   x"15", 
  x"73",   x"79",   x"67",   x"6D",   x"5B",   x"51",   x"4F",   x"45", 
  x"C5",   x"CF",   x"D1",   x"DB",   x"ED",   x"E7",   x"F9",   x"F3", 
  x"95",   x"9F",   x"81",   x"8B",   x"BD",   x"B7",   x"A9",   x"A3", 
  x"65",   x"6F",   x"71",   x"7B",   x"4D",   x"47",   x"59",   x"53", 
  x"35",   x"3F",   x"21",   x"2B",   x"1D",   x"17",   x"09",   x"03", 
  x"46",   x"4C",   x"52",   x"58",   x"6E",   x"64",   x"7A",   x"70", 
  x"16",   x"1C",   x"02",   x"08",   x"3E",   x"34",   x"2A",   x"20", 
  x"E6",   x"EC",   x"F2",   x"F8",   x"CE",   x"C4",   x"DA",   x"D0", 
  x"B6",   x"BC",   x"A2",   x"A8",   x"9E",   x"94",   x"8A",   x"80", 
  x"49",   x"43",   x"5D",   x"57",   x"61",   x"6B",   x"75",   x"7F", 
  x"19",   x"13",   x"0D",   x"07",   x"31",   x"3B",   x"25",   x"2F", 
  x"E9",   x"E3",   x"FD",   x"F7",   x"C1",   x"CB",   x"D5",   x"DF", 
  x"B9",   x"B3",   x"AD",   x"A7",   x"91",   x"9B",   x"85",   x"8F", 
  x"CA",   x"C0",   x"DE",   x"D4",   x"E2",   x"E8",   x"F6",   x"FC", 
  x"9A",   x"90",   x"8E",   x"84",   x"B2",   x"B8",   x"A6",   x"AC", 
  x"6A",   x"60",   x"7E",   x"74",   x"42",   x"48",   x"56",   x"5C", 
  x"3A",   x"30",   x"2E",   x"24",   x"12",   x"18",   x"06",   x"0C", 
  x"8C",   x"86",   x"98",   x"92",   x"A4",   x"AE",   x"B0",   x"BA", 
  x"DC",   x"D6",   x"C8",   x"C2",   x"F4",   x"FE",   x"E0",   x"EA", 
  x"2C",   x"26",   x"38",   x"32",   x"04",   x"0E",   x"10",   x"1A", 
  x"7C",   x"76",   x"68",   x"62",   x"54",   x"5E",   x"40",   x"4A", 
  x"0F",   x"05",   x"1B",   x"11",   x"27",   x"2D",   x"33",   x"39", 
  x"5F",   x"55",   x"4B",   x"41",   x"77",   x"7D",   x"63",   x"69", 
  x"AF",   x"A5",   x"BB",   x"B1",   x"87",   x"8D",   x"93",   x"99", 
  x"FF",   x"F5",   x"EB",   x"E1",   x"D7",   x"DD",   x"C3",   x"C9", 
  x"00",   x"0B",   x"16",   x"1D",   x"2C",   x"27",   x"3A",   x"31", 
  x"58",   x"53",   x"4E",   x"45",   x"74",   x"7F",   x"62",   x"69", 
  x"B0",   x"BB",   x"A6",   x"AD",   x"9C",   x"97",   x"8A",   x"81", 
  x"E8",   x"E3",   x"FE",   x"F5",   x"C4",   x"CF",   x"D2",   x"D9", 
  x"A3",   x"A8",   x"B5",   x"BE",   x"8F",   x"84",   x"99",   x"92", 
  x"FB",   x"F0",   x"ED",   x"E6",   x"D7",   x"DC",   x"C1",   x"CA", 
  x"13",   x"18",   x"05",   x"0E",   x"3F",   x"34",   x"29",   x"22", 
  x"4B",   x"40",   x"5D",   x"56",   x"67",   x"6C",   x"71",   x"7A", 
  x"85",   x"8E",   x"93",   x"98",   x"A9",   x"A2",   x"BF",   x"B4", 
  x"DD",   x"D6",   x"CB",   x"C0",   x"F1",   x"FA",   x"E7",   x"EC", 
  x"35",   x"3E",   x"23",   x"28",   x"19",   x"12",   x"0F",   x"04", 
  x"6D",   x"66",   x"7B",   x"70",   x"41",   x"4A",   x"57",   x"5C", 
  x"26",   x"2D",   x"30",   x"3B",   x"0A",   x"01",   x"1C",   x"17", 
  x"7E",   x"75",   x"68",   x"63",   x"52",   x"59",   x"44",   x"4F", 
  x"96",   x"9D",   x"80",   x"8B",   x"BA",   x"B1",   x"AC",   x"A7", 
  x"CE",   x"C5",   x"D8",   x"D3",   x"E2",   x"E9",   x"F4",   x"FF", 
  x"C9",   x"C2",   x"DF",   x"D4",   x"E5",   x"EE",   x"F3",   x"F8", 
  x"91",   x"9A",   x"87",   x"8C",   x"BD",   x"B6",   x"AB",   x"A0", 
  x"79",   x"72",   x"6F",   x"64",   x"55",   x"5E",   x"43",   x"48", 
  x"21",   x"2A",   x"37",   x"3C",   x"0D",   x"06",   x"1B",   x"10", 
  x"6A",   x"61",   x"7C",   x"77",   x"46",   x"4D",   x"50",   x"5B", 
  x"32",   x"39",   x"24",   x"2F",   x"1E",   x"15",   x"08",   x"03", 
  x"DA",   x"D1",   x"CC",   x"C7",   x"F6",   x"FD",   x"E0",   x"EB", 
  x"82",   x"89",   x"94",   x"9F",   x"AE",   x"A5",   x"B8",   x"B3", 
  x"4C",   x"47",   x"5A",   x"51",   x"60",   x"6B",   x"76",   x"7D", 
  x"14",   x"1F",   x"02",   x"09",   x"38",   x"33",   x"2E",   x"25", 
  x"FC",   x"F7",   x"EA",   x"E1",   x"D0",   x"DB",   x"C6",   x"CD", 
  x"A4",   x"AF",   x"B2",   x"B9",   x"88",   x"83",   x"9E",   x"95", 
  x"EF",   x"E4",   x"F9",   x"F2",   x"C3",   x"C8",   x"D5",   x"DE", 
  x"B7",   x"BC",   x"A1",   x"AA",   x"9B",   x"90",   x"8D",   x"86", 
  x"5F",   x"54",   x"49",   x"42",   x"73",   x"78",   x"65",   x"6E", 
  x"07",   x"0C",   x"11",   x"1A",   x"2B",   x"20",   x"3D",   x"36", 
  x"00",   x"0C",   x"18",   x"14",   x"30",   x"3C",   x"28",   x"24", 
  x"60",   x"6C",   x"78",   x"74",   x"50",   x"5C",   x"48",   x"44", 
  x"C0",   x"CC",   x"D8",   x"D4",   x"F0",   x"FC",   x"E8",   x"E4", 
  x"A0",   x"AC",   x"B8",   x"B4",   x"90",   x"9C",   x"88",   x"84", 
  x"43",   x"4F",   x"5B",   x"57",   x"73",   x"7F",   x"6B",   x"67", 
  x"23",   x"2F",   x"3B",   x"37",   x"13",   x"1F",   x"0B",   x"07", 
  x"83",   x"8F",   x"9B",   x"97",   x"B3",   x"BF",   x"AB",   x"A7", 
  x"E3",   x"EF",   x"FB",   x"F7",   x"D3",   x"DF",   x"CB",   x"C7", 
  x"86",   x"8A",   x"9E",   x"92",   x"B6",   x"BA",   x"AE",   x"A2", 
  x"E6",   x"EA",   x"FE",   x"F2",   x"D6",   x"DA",   x"CE",   x"C2", 
  x"46",   x"4A",   x"5E",   x"52",   x"76",   x"7A",   x"6E",   x"62", 
  x"26",   x"2A",   x"3E",   x"32",   x"16",   x"1A",   x"0E",   x"02", 
  x"C5",   x"C9",   x"DD",   x"D1",   x"F5",   x"F9",   x"ED",   x"E1", 
  x"A5",   x"A9",   x"BD",   x"B1",   x"95",   x"99",   x"8D",   x"81", 
  x"05",   x"09",   x"1D",   x"11",   x"35",   x"39",   x"2D",   x"21", 
  x"65",   x"69",   x"7D",   x"71",   x"55",   x"59",   x"4D",   x"41", 
  x"CF",   x"C3",   x"D7",   x"DB",   x"FF",   x"F3",   x"E7",   x"EB", 
  x"AF",   x"A3",   x"B7",   x"BB",   x"9F",   x"93",   x"87",   x"8B", 
  x"0F",   x"03",   x"17",   x"1B",   x"3F",   x"33",   x"27",   x"2B", 
  x"6F",   x"63",   x"77",   x"7B",   x"5F",   x"53",   x"47",   x"4B", 
  x"8C",   x"80",   x"94",   x"98",   x"BC",   x"B0",   x"A4",   x"A8", 
  x"EC",   x"E0",   x"F4",   x"F8",   x"DC",   x"D0",   x"C4",   x"C8", 
  x"4C",   x"40",   x"54",   x"58",   x"7C",   x"70",   x"64",   x"68", 
  x"2C",   x"20",   x"34",   x"38",   x"1C",   x"10",   x"04",   x"08", 
  x"49",   x"45",   x"51",   x"5D",   x"79",   x"75",   x"61",   x"6D", 
  x"29",   x"25",   x"31",   x"3D",   x"19",   x"15",   x"01",   x"0D", 
  x"89",   x"85",   x"91",   x"9D",   x"B9",   x"B5",   x"A1",   x"AD", 
  x"E9",   x"E5",   x"F1",   x"FD",   x"D9",   x"D5",   x"C1",   x"CD", 
  x"0A",   x"06",   x"12",   x"1E",   x"3A",   x"36",   x"22",   x"2E", 
  x"6A",   x"66",   x"72",   x"7E",   x"5A",   x"56",   x"42",   x"4E", 
  x"CA",   x"C6",   x"D2",   x"DE",   x"FA",   x"F6",   x"E2",   x"EE", 
  x"AA",   x"A6",   x"B2",   x"BE",   x"9A",   x"96",   x"82",   x"8E", 
  x"00",   x"0D",   x"1A",   x"17",   x"34",   x"39",   x"2E",   x"23", 
  x"68",   x"65",   x"72",   x"7F",   x"5C",   x"51",   x"46",   x"4B", 
  x"D0",   x"DD",   x"CA",   x"C7",   x"E4",   x"E9",   x"FE",   x"F3", 
  x"B8",   x"B5",   x"A2",   x"AF",   x"8C",   x"81",   x"96",   x"9B", 
  x"63",   x"6E",   x"79",   x"74",   x"57",   x"5A",   x"4D",   x"40", 
  x"0B",   x"06",   x"11",   x"1C",   x"3F",   x"32",   x"25",   x"28", 
  x"B3",   x"BE",   x"A9",   x"A4",   x"87",   x"8A",   x"9D",   x"90", 
  x"DB",   x"D6",   x"C1",   x"CC",   x"EF",   x"E2",   x"F5",   x"F8", 
  x"C6",   x"CB",   x"DC",   x"D1",   x"F2",   x"FF",   x"E8",   x"E5", 
  x"AE",   x"A3",   x"B4",   x"B9",   x"9A",   x"97",   x"80",   x"8D", 
  x"16",   x"1B",   x"0C",   x"01",   x"22",   x"2F",   x"38",   x"35", 
  x"7E",   x"73",   x"64",   x"69",   x"4A",   x"47",   x"50",   x"5D", 
  x"A5",   x"A8",   x"BF",   x"B2",   x"91",   x"9C",   x"8B",   x"86", 
  x"CD",   x"C0",   x"D7",   x"DA",   x"F9",   x"F4",   x"E3",   x"EE", 
  x"75",   x"78",   x"6F",   x"62",   x"41",   x"4C",   x"5B",   x"56", 
  x"1D",   x"10",   x"07",   x"0A",   x"29",   x"24",   x"33",   x"3E", 
  x"4F",   x"42",   x"55",   x"58",   x"7B",   x"76",   x"61",   x"6C", 
  x"27",   x"2A",   x"3D",   x"30",   x"13",   x"1E",   x"09",   x"04", 
  x"9F",   x"92",   x"85",   x"88",   x"AB",   x"A6",   x"B1",   x"BC", 
  x"F7",   x"FA",   x"ED",   x"E0",   x"C3",   x"CE",   x"D9",   x"D4", 
  x"2C",   x"21",   x"36",   x"3B",   x"18",   x"15",   x"02",   x"0F", 
  x"44",   x"49",   x"5E",   x"53",   x"70",   x"7D",   x"6A",   x"67", 
  x"FC",   x"F1",   x"E6",   x"EB",   x"C8",   x"C5",   x"D2",   x"DF", 
  x"94",   x"99",   x"8E",   x"83",   x"A0",   x"AD",   x"BA",   x"B7", 
  x"89",   x"84",   x"93",   x"9E",   x"BD",   x"B0",   x"A7",   x"AA", 
  x"E1",   x"EC",   x"FB",   x"F6",   x"D5",   x"D8",   x"CF",   x"C2", 
  x"59",   x"54",   x"43",   x"4E",   x"6D",   x"60",   x"77",   x"7A", 
  x"31",   x"3C",   x"2B",   x"26",   x"05",   x"08",   x"1F",   x"12", 
  x"EA",   x"E7",   x"F0",   x"FD",   x"DE",   x"D3",   x"C4",   x"C9", 
  x"82",   x"8F",   x"98",   x"95",   x"B6",   x"BB",   x"AC",   x"A1", 
  x"3A",   x"37",   x"20",   x"2D",   x"0E",   x"03",   x"14",   x"19", 
  x"52",   x"5F",   x"48",   x"45",   x"66",   x"6B",   x"7C",   x"71", 
  x"00",   x"0E",   x"1C",   x"12",   x"38",   x"36",   x"24",   x"2A", 
  x"70",   x"7E",   x"6C",   x"62",   x"48",   x"46",   x"54",   x"5A", 
  x"E0",   x"EE",   x"FC",   x"F2",   x"D8",   x"D6",   x"C4",   x"CA", 
  x"90",   x"9E",   x"8C",   x"82",   x"A8",   x"A6",   x"B4",   x"BA", 
  x"03",   x"0D",   x"1F",   x"11",   x"3B",   x"35",   x"27",   x"29", 
  x"73",   x"7D",   x"6F",   x"61",   x"4B",   x"45",   x"57",   x"59", 
  x"E3",   x"ED",   x"FF",   x"F1",   x"DB",   x"D5",   x"C7",   x"C9", 
  x"93",   x"9D",   x"8F",   x"81",   x"AB",   x"A5",   x"B7",   x"B9", 
  x"06",   x"08",   x"1A",   x"14",   x"3E",   x"30",   x"22",   x"2C", 
  x"76",   x"78",   x"6A",   x"64",   x"4E",   x"40",   x"52",   x"5C", 
  x"E6",   x"E8",   x"FA",   x"F4",   x"DE",   x"D0",   x"C2",   x"CC", 
  x"96",   x"98",   x"8A",   x"84",   x"AE",   x"A0",   x"B2",   x"BC", 
  x"05",   x"0B",   x"19",   x"17",   x"3D",   x"33",   x"21",   x"2F", 
  x"75",   x"7B",   x"69",   x"67",   x"4D",   x"43",   x"51",   x"5F", 
  x"E5",   x"EB",   x"F9",   x"F7",   x"DD",   x"D3",   x"C1",   x"CF", 
  x"95",   x"9B",   x"89",   x"87",   x"AD",   x"A3",   x"B1",   x"BF", 
  x"0C",   x"02",   x"10",   x"1E",   x"34",   x"3A",   x"28",   x"26", 
  x"7C",   x"72",   x"60",   x"6E",   x"44",   x"4A",   x"58",   x"56", 
  x"EC",   x"E2",   x"F0",   x"FE",   x"D4",   x"DA",   x"C8",   x"C6", 
  x"9C",   x"92",   x"80",   x"8E",   x"A4",   x"AA",   x"B8",   x"B6", 
  x"0F",   x"01",   x"13",   x"1D",   x"37",   x"39",   x"2B",   x"25", 
  x"7F",   x"71",   x"63",   x"6D",   x"47",   x"49",   x"5B",   x"55", 
  x"EF",   x"E1",   x"F3",   x"FD",   x"D7",   x"D9",   x"CB",   x"C5", 
  x"9F",   x"91",   x"83",   x"8D",   x"A7",   x"A9",   x"BB",   x"B5", 
  x"0A",   x"04",   x"16",   x"18",   x"32",   x"3C",   x"2E",   x"20", 
  x"7A",   x"74",   x"66",   x"68",   x"42",   x"4C",   x"5E",   x"50", 
  x"EA",   x"E4",   x"F6",   x"F8",   x"D2",   x"DC",   x"CE",   x"C0", 
  x"9A",   x"94",   x"86",   x"88",   x"A2",   x"AC",   x"BE",   x"B0", 
  x"09",   x"07",   x"15",   x"1B",   x"31",   x"3F",   x"2D",   x"23", 
  x"79",   x"77",   x"65",   x"6B",   x"41",   x"4F",   x"5D",   x"53", 
  x"E9",   x"E7",   x"F5",   x"FB",   x"D1",   x"DF",   x"CD",   x"C3", 
  x"99",   x"97",   x"85",   x"8B",   x"A1",   x"AF",   x"BD",   x"B3", 
  x"00",   x"0F",   x"1E",   x"11",   x"3C",   x"33",   x"22",   x"2D", 
  x"78",   x"77",   x"66",   x"69",   x"44",   x"4B",   x"5A",   x"55", 
  x"F0",   x"FF",   x"EE",   x"E1",   x"CC",   x"C3",   x"D2",   x"DD", 
  x"88",   x"87",   x"96",   x"99",   x"B4",   x"BB",   x"AA",   x"A5", 
  x"23",   x"2C",   x"3D",   x"32",   x"1F",   x"10",   x"01",   x"0E", 
  x"5B",   x"54",   x"45",   x"4A",   x"67",   x"68",   x"79",   x"76", 
  x"D3",   x"DC",   x"CD",   x"C2",   x"EF",   x"E0",   x"F1",   x"FE", 
  x"AB",   x"A4",   x"B5",   x"BA",   x"97",   x"98",   x"89",   x"86", 
  x"46",   x"49",   x"58",   x"57",   x"7A",   x"75",   x"64",   x"6B", 
  x"3E",   x"31",   x"20",   x"2F",   x"02",   x"0D",   x"1C",   x"13", 
  x"B6",   x"B9",   x"A8",   x"A7",   x"8A",   x"85",   x"94",   x"9B", 
  x"CE",   x"C1",   x"D0",   x"DF",   x"F2",   x"FD",   x"EC",   x"E3", 
  x"65",   x"6A",   x"7B",   x"74",   x"59",   x"56",   x"47",   x"48", 
  x"1D",   x"12",   x"03",   x"0C",   x"21",   x"2E",   x"3F",   x"30", 
  x"95",   x"9A",   x"8B",   x"84",   x"A9",   x"A6",   x"B7",   x"B8", 
  x"ED",   x"E2",   x"F3",   x"FC",   x"D1",   x"DE",   x"CF",   x"C0", 
  x"8C",   x"83",   x"92",   x"9D",   x"B0",   x"BF",   x"AE",   x"A1", 
  x"F4",   x"FB",   x"EA",   x"E5",   x"C8",   x"C7",   x"D6",   x"D9", 
  x"7C",   x"73",   x"62",   x"6D",   x"40",   x"4F",   x"5E",   x"51", 
  x"04",   x"0B",   x"1A",   x"15",   x"38",   x"37",   x"26",   x"29", 
  x"AF",   x"A0",   x"B1",   x"BE",   x"93",   x"9C",   x"8D",   x"82", 
  x"D7",   x"D8",   x"C9",   x"C6",   x"EB",   x"E4",   x"F5",   x"FA", 
  x"5F",   x"50",   x"41",   x"4E",   x"63",   x"6C",   x"7D",   x"72", 
  x"27",   x"28",   x"39",   x"36",   x"1B",   x"14",   x"05",   x"0A", 
  x"CA",   x"C5",   x"D4",   x"DB",   x"F6",   x"F9",   x"E8",   x"E7", 
  x"B2",   x"BD",   x"AC",   x"A3",   x"8E",   x"81",   x"90",   x"9F", 
  x"3A",   x"35",   x"24",   x"2B",   x"06",   x"09",   x"18",   x"17", 
  x"42",   x"4D",   x"5C",   x"53",   x"7E",   x"71",   x"60",   x"6F", 
  x"E9",   x"E6",   x"F7",   x"F8",   x"D5",   x"DA",   x"CB",   x"C4", 
  x"91",   x"9E",   x"8F",   x"80",   x"AD",   x"A2",   x"B3",   x"BC", 
  x"19",   x"16",   x"07",   x"08",   x"25",   x"2A",   x"3B",   x"34", 
  x"61",   x"6E",   x"7F",   x"70",   x"5D",   x"52",   x"43",   x"4C", 
  x"00",   x"10",   x"20",   x"30",   x"40",   x"50",   x"60",   x"70", 
  x"80",   x"90",   x"A0",   x"B0",   x"C0",   x"D0",   x"E0",   x"F0", 
  x"C3",   x"D3",   x"E3",   x"F3",   x"83",   x"93",   x"A3",   x"B3", 
  x"43",   x"53",   x"63",   x"73",   x"03",   x"13",   x"23",   x"33", 
  x"45",   x"55",   x"65",   x"75",   x"05",   x"15",   x"25",   x"35", 
  x"C5",   x"D5",   x"E5",   x"F5",   x"85",   x"95",   x"A5",   x"B5", 
  x"86",   x"96",   x"A6",   x"B6",   x"C6",   x"D6",   x"E6",   x"F6", 
  x"06",   x"16",   x"26",   x"36",   x"46",   x"56",   x"66",   x"76", 
  x"8A",   x"9A",   x"AA",   x"BA",   x"CA",   x"DA",   x"EA",   x"FA", 
  x"0A",   x"1A",   x"2A",   x"3A",   x"4A",   x"5A",   x"6A",   x"7A", 
  x"49",   x"59",   x"69",   x"79",   x"09",   x"19",   x"29",   x"39", 
  x"C9",   x"D9",   x"E9",   x"F9",   x"89",   x"99",   x"A9",   x"B9", 
  x"CF",   x"DF",   x"EF",   x"FF",   x"8F",   x"9F",   x"AF",   x"BF", 
  x"4F",   x"5F",   x"6F",   x"7F",   x"0F",   x"1F",   x"2F",   x"3F", 
  x"0C",   x"1C",   x"2C",   x"3C",   x"4C",   x"5C",   x"6C",   x"7C", 
  x"8C",   x"9C",   x"AC",   x"BC",   x"CC",   x"DC",   x"EC",   x"FC", 
  x"D7",   x"C7",   x"F7",   x"E7",   x"97",   x"87",   x"B7",   x"A7", 
  x"57",   x"47",   x"77",   x"67",   x"17",   x"07",   x"37",   x"27", 
  x"14",   x"04",   x"34",   x"24",   x"54",   x"44",   x"74",   x"64", 
  x"94",   x"84",   x"B4",   x"A4",   x"D4",   x"C4",   x"F4",   x"E4", 
  x"92",   x"82",   x"B2",   x"A2",   x"D2",   x"C2",   x"F2",   x"E2", 
  x"12",   x"02",   x"32",   x"22",   x"52",   x"42",   x"72",   x"62", 
  x"51",   x"41",   x"71",   x"61",   x"11",   x"01",   x"31",   x"21", 
  x"D1",   x"C1",   x"F1",   x"E1",   x"91",   x"81",   x"B1",   x"A1", 
  x"5D",   x"4D",   x"7D",   x"6D",   x"1D",   x"0D",   x"3D",   x"2D", 
  x"DD",   x"CD",   x"FD",   x"ED",   x"9D",   x"8D",   x"BD",   x"AD", 
  x"9E",   x"8E",   x"BE",   x"AE",   x"DE",   x"CE",   x"FE",   x"EE", 
  x"1E",   x"0E",   x"3E",   x"2E",   x"5E",   x"4E",   x"7E",   x"6E", 
  x"18",   x"08",   x"38",   x"28",   x"58",   x"48",   x"78",   x"68", 
  x"98",   x"88",   x"B8",   x"A8",   x"D8",   x"C8",   x"F8",   x"E8", 
  x"DB",   x"CB",   x"FB",   x"EB",   x"9B",   x"8B",   x"BB",   x"AB", 
  x"5B",   x"4B",   x"7B",   x"6B",   x"1B",   x"0B",   x"3B",   x"2B", 
  x"00",   x"11",   x"22",   x"33",   x"44",   x"55",   x"66",   x"77", 
  x"88",   x"99",   x"AA",   x"BB",   x"CC",   x"DD",   x"EE",   x"FF", 
  x"D3",   x"C2",   x"F1",   x"E0",   x"97",   x"86",   x"B5",   x"A4", 
  x"5B",   x"4A",   x"79",   x"68",   x"1F",   x"0E",   x"3D",   x"2C", 
  x"65",   x"74",   x"47",   x"56",   x"21",   x"30",   x"03",   x"12", 
  x"ED",   x"FC",   x"CF",   x"DE",   x"A9",   x"B8",   x"8B",   x"9A", 
  x"B6",   x"A7",   x"94",   x"85",   x"F2",   x"E3",   x"D0",   x"C1", 
  x"3E",   x"2F",   x"1C",   x"0D",   x"7A",   x"6B",   x"58",   x"49", 
  x"CA",   x"DB",   x"E8",   x"F9",   x"8E",   x"9F",   x"AC",   x"BD", 
  x"42",   x"53",   x"60",   x"71",   x"06",   x"17",   x"24",   x"35", 
  x"19",   x"08",   x"3B",   x"2A",   x"5D",   x"4C",   x"7F",   x"6E", 
  x"91",   x"80",   x"B3",   x"A2",   x"D5",   x"C4",   x"F7",   x"E6", 
  x"AF",   x"BE",   x"8D",   x"9C",   x"EB",   x"FA",   x"C9",   x"D8", 
  x"27",   x"36",   x"05",   x"14",   x"63",   x"72",   x"41",   x"50", 
  x"7C",   x"6D",   x"5E",   x"4F",   x"38",   x"29",   x"1A",   x"0B", 
  x"F4",   x"E5",   x"D6",   x"C7",   x"B0",   x"A1",   x"92",   x"83", 
  x"57",   x"46",   x"75",   x"64",   x"13",   x"02",   x"31",   x"20", 
  x"DF",   x"CE",   x"FD",   x"EC",   x"9B",   x"8A",   x"B9",   x"A8", 
  x"84",   x"95",   x"A6",   x"B7",   x"C0",   x"D1",   x"E2",   x"F3", 
  x"0C",   x"1D",   x"2E",   x"3F",   x"48",   x"59",   x"6A",   x"7B", 
  x"32",   x"23",   x"10",   x"01",   x"76",   x"67",   x"54",   x"45", 
  x"BA",   x"AB",   x"98",   x"89",   x"FE",   x"EF",   x"DC",   x"CD", 
  x"E1",   x"F0",   x"C3",   x"D2",   x"A5",   x"B4",   x"87",   x"96", 
  x"69",   x"78",   x"4B",   x"5A",   x"2D",   x"3C",   x"0F",   x"1E", 
  x"9D",   x"8C",   x"BF",   x"AE",   x"D9",   x"C8",   x"FB",   x"EA", 
  x"15",   x"04",   x"37",   x"26",   x"51",   x"40",   x"73",   x"62", 
  x"4E",   x"5F",   x"6C",   x"7D",   x"0A",   x"1B",   x"28",   x"39", 
  x"C6",   x"D7",   x"E4",   x"F5",   x"82",   x"93",   x"A0",   x"B1", 
  x"F8",   x"E9",   x"DA",   x"CB",   x"BC",   x"AD",   x"9E",   x"8F", 
  x"70",   x"61",   x"52",   x"43",   x"34",   x"25",   x"16",   x"07", 
  x"2B",   x"3A",   x"09",   x"18",   x"6F",   x"7E",   x"4D",   x"5C", 
  x"A3",   x"B2",   x"81",   x"90",   x"E7",   x"F6",   x"C5",   x"D4", 
  x"00",   x"12",   x"24",   x"36",   x"48",   x"5A",   x"6C",   x"7E", 
  x"90",   x"82",   x"B4",   x"A6",   x"D8",   x"CA",   x"FC",   x"EE", 
  x"E3",   x"F1",   x"C7",   x"D5",   x"AB",   x"B9",   x"8F",   x"9D", 
  x"73",   x"61",   x"57",   x"45",   x"3B",   x"29",   x"1F",   x"0D", 
  x"05",   x"17",   x"21",   x"33",   x"4D",   x"5F",   x"69",   x"7B", 
  x"95",   x"87",   x"B1",   x"A3",   x"DD",   x"CF",   x"F9",   x"EB", 
  x"E6",   x"F4",   x"C2",   x"D0",   x"AE",   x"BC",   x"8A",   x"98", 
  x"76",   x"64",   x"52",   x"40",   x"3E",   x"2C",   x"1A",   x"08", 
  x"0A",   x"18",   x"2E",   x"3C",   x"42",   x"50",   x"66",   x"74", 
  x"9A",   x"88",   x"BE",   x"AC",   x"D2",   x"C0",   x"F6",   x"E4", 
  x"E9",   x"FB",   x"CD",   x"DF",   x"A1",   x"B3",   x"85",   x"97", 
  x"79",   x"6B",   x"5D",   x"4F",   x"31",   x"23",   x"15",   x"07", 
  x"0F",   x"1D",   x"2B",   x"39",   x"47",   x"55",   x"63",   x"71", 
  x"9F",   x"8D",   x"BB",   x"A9",   x"D7",   x"C5",   x"F3",   x"E1", 
  x"EC",   x"FE",   x"C8",   x"DA",   x"A4",   x"B6",   x"80",   x"92", 
  x"7C",   x"6E",   x"58",   x"4A",   x"34",   x"26",   x"10",   x"02", 
  x"14",   x"06",   x"30",   x"22",   x"5C",   x"4E",   x"78",   x"6A", 
  x"84",   x"96",   x"A0",   x"B2",   x"CC",   x"DE",   x"E8",   x"FA", 
  x"F7",   x"E5",   x"D3",   x"C1",   x"BF",   x"AD",   x"9B",   x"89", 
  x"67",   x"75",   x"43",   x"51",   x"2F",   x"3D",   x"0B",   x"19", 
  x"11",   x"03",   x"35",   x"27",   x"59",   x"4B",   x"7D",   x"6F", 
  x"81",   x"93",   x"A5",   x"B7",   x"C9",   x"DB",   x"ED",   x"FF", 
  x"F2",   x"E0",   x"D6",   x"C4",   x"BA",   x"A8",   x"9E",   x"8C", 
  x"62",   x"70",   x"46",   x"54",   x"2A",   x"38",   x"0E",   x"1C", 
  x"1E",   x"0C",   x"3A",   x"28",   x"56",   x"44",   x"72",   x"60", 
  x"8E",   x"9C",   x"AA",   x"B8",   x"C6",   x"D4",   x"E2",   x"F0", 
  x"FD",   x"EF",   x"D9",   x"CB",   x"B5",   x"A7",   x"91",   x"83", 
  x"6D",   x"7F",   x"49",   x"5B",   x"25",   x"37",   x"01",   x"13", 
  x"1B",   x"09",   x"3F",   x"2D",   x"53",   x"41",   x"77",   x"65", 
  x"8B",   x"99",   x"AF",   x"BD",   x"C3",   x"D1",   x"E7",   x"F5", 
  x"F8",   x"EA",   x"DC",   x"CE",   x"B0",   x"A2",   x"94",   x"86", 
  x"68",   x"7A",   x"4C",   x"5E",   x"20",   x"32",   x"04",   x"16", 
  x"00",   x"13",   x"26",   x"35",   x"4C",   x"5F",   x"6A",   x"79", 
  x"98",   x"8B",   x"BE",   x"AD",   x"D4",   x"C7",   x"F2",   x"E1", 
  x"F3",   x"E0",   x"D5",   x"C6",   x"BF",   x"AC",   x"99",   x"8A", 
  x"6B",   x"78",   x"4D",   x"5E",   x"27",   x"34",   x"01",   x"12", 
  x"25",   x"36",   x"03",   x"10",   x"69",   x"7A",   x"4F",   x"5C", 
  x"BD",   x"AE",   x"9B",   x"88",   x"F1",   x"E2",   x"D7",   x"C4", 
  x"D6",   x"C5",   x"F0",   x"E3",   x"9A",   x"89",   x"BC",   x"AF", 
  x"4E",   x"5D",   x"68",   x"7B",   x"02",   x"11",   x"24",   x"37", 
  x"4A",   x"59",   x"6C",   x"7F",   x"06",   x"15",   x"20",   x"33", 
  x"D2",   x"C1",   x"F4",   x"E7",   x"9E",   x"8D",   x"B8",   x"AB", 
  x"B9",   x"AA",   x"9F",   x"8C",   x"F5",   x"E6",   x"D3",   x"C0", 
  x"21",   x"32",   x"07",   x"14",   x"6D",   x"7E",   x"4B",   x"58", 
  x"6F",   x"7C",   x"49",   x"5A",   x"23",   x"30",   x"05",   x"16", 
  x"F7",   x"E4",   x"D1",   x"C2",   x"BB",   x"A8",   x"9D",   x"8E", 
  x"9C",   x"8F",   x"BA",   x"A9",   x"D0",   x"C3",   x"F6",   x"E5", 
  x"04",   x"17",   x"22",   x"31",   x"48",   x"5B",   x"6E",   x"7D", 
  x"94",   x"87",   x"B2",   x"A1",   x"D8",   x"CB",   x"FE",   x"ED", 
  x"0C",   x"1F",   x"2A",   x"39",   x"40",   x"53",   x"66",   x"75", 
  x"67",   x"74",   x"41",   x"52",   x"2B",   x"38",   x"0D",   x"1E", 
  x"FF",   x"EC",   x"D9",   x"CA",   x"B3",   x"A0",   x"95",   x"86", 
  x"B1",   x"A2",   x"97",   x"84",   x"FD",   x"EE",   x"DB",   x"C8", 
  x"29",   x"3A",   x"0F",   x"1C",   x"65",   x"76",   x"43",   x"50", 
  x"42",   x"51",   x"64",   x"77",   x"0E",   x"1D",   x"28",   x"3B", 
  x"DA",   x"C9",   x"FC",   x"EF",   x"96",   x"85",   x"B0",   x"A3", 
  x"DE",   x"CD",   x"F8",   x"EB",   x"92",   x"81",   x"B4",   x"A7", 
  x"46",   x"55",   x"60",   x"73",   x"0A",   x"19",   x"2C",   x"3F", 
  x"2D",   x"3E",   x"0B",   x"18",   x"61",   x"72",   x"47",   x"54", 
  x"B5",   x"A6",   x"93",   x"80",   x"F9",   x"EA",   x"DF",   x"CC", 
  x"FB",   x"E8",   x"DD",   x"CE",   x"B7",   x"A4",   x"91",   x"82", 
  x"63",   x"70",   x"45",   x"56",   x"2F",   x"3C",   x"09",   x"1A", 
  x"08",   x"1B",   x"2E",   x"3D",   x"44",   x"57",   x"62",   x"71", 
  x"90",   x"83",   x"B6",   x"A5",   x"DC",   x"CF",   x"FA",   x"E9", 
  x"00",   x"14",   x"28",   x"3C",   x"50",   x"44",   x"78",   x"6C", 
  x"A0",   x"B4",   x"88",   x"9C",   x"F0",   x"E4",   x"D8",   x"CC", 
  x"83",   x"97",   x"AB",   x"BF",   x"D3",   x"C7",   x"FB",   x"EF", 
  x"23",   x"37",   x"0B",   x"1F",   x"73",   x"67",   x"5B",   x"4F", 
  x"C5",   x"D1",   x"ED",   x"F9",   x"95",   x"81",   x"BD",   x"A9", 
  x"65",   x"71",   x"4D",   x"59",   x"35",   x"21",   x"1D",   x"09", 
  x"46",   x"52",   x"6E",   x"7A",   x"16",   x"02",   x"3E",   x"2A", 
  x"E6",   x"F2",   x"CE",   x"DA",   x"B6",   x"A2",   x"9E",   x"8A", 
  x"49",   x"5D",   x"61",   x"75",   x"19",   x"0D",   x"31",   x"25", 
  x"E9",   x"FD",   x"C1",   x"D5",   x"B9",   x"AD",   x"91",   x"85", 
  x"CA",   x"DE",   x"E2",   x"F6",   x"9A",   x"8E",   x"B2",   x"A6", 
  x"6A",   x"7E",   x"42",   x"56",   x"3A",   x"2E",   x"12",   x"06", 
  x"8C",   x"98",   x"A4",   x"B0",   x"DC",   x"C8",   x"F4",   x"E0", 
  x"2C",   x"38",   x"04",   x"10",   x"7C",   x"68",   x"54",   x"40", 
  x"0F",   x"1B",   x"27",   x"33",   x"5F",   x"4B",   x"77",   x"63", 
  x"AF",   x"BB",   x"87",   x"93",   x"FF",   x"EB",   x"D7",   x"C3", 
  x"92",   x"86",   x"BA",   x"AE",   x"C2",   x"D6",   x"EA",   x"FE", 
  x"32",   x"26",   x"1A",   x"0E",   x"62",   x"76",   x"4A",   x"5E", 
  x"11",   x"05",   x"39",   x"2D",   x"41",   x"55",   x"69",   x"7D", 
  x"B1",   x"A5",   x"99",   x"8D",   x"E1",   x"F5",   x"C9",   x"DD", 
  x"57",   x"43",   x"7F",   x"6B",   x"07",   x"13",   x"2F",   x"3B", 
  x"F7",   x"E3",   x"DF",   x"CB",   x"A7",   x"B3",   x"8F",   x"9B", 
  x"D4",   x"C0",   x"FC",   x"E8",   x"84",   x"90",   x"AC",   x"B8", 
  x"74",   x"60",   x"5C",   x"48",   x"24",   x"30",   x"0C",   x"18", 
  x"DB",   x"CF",   x"F3",   x"E7",   x"8B",   x"9F",   x"A3",   x"B7", 
  x"7B",   x"6F",   x"53",   x"47",   x"2B",   x"3F",   x"03",   x"17", 
  x"58",   x"4C",   x"70",   x"64",   x"08",   x"1C",   x"20",   x"34", 
  x"F8",   x"EC",   x"D0",   x"C4",   x"A8",   x"BC",   x"80",   x"94", 
  x"1E",   x"0A",   x"36",   x"22",   x"4E",   x"5A",   x"66",   x"72", 
  x"BE",   x"AA",   x"96",   x"82",   x"EE",   x"FA",   x"C6",   x"D2", 
  x"9D",   x"89",   x"B5",   x"A1",   x"CD",   x"D9",   x"E5",   x"F1", 
  x"3D",   x"29",   x"15",   x"01",   x"6D",   x"79",   x"45",   x"51", 
  x"00",   x"15",   x"2A",   x"3F",   x"54",   x"41",   x"7E",   x"6B", 
  x"A8",   x"BD",   x"82",   x"97",   x"FC",   x"E9",   x"D6",   x"C3", 
  x"93",   x"86",   x"B9",   x"AC",   x"C7",   x"D2",   x"ED",   x"F8", 
  x"3B",   x"2E",   x"11",   x"04",   x"6F",   x"7A",   x"45",   x"50", 
  x"E5",   x"F0",   x"CF",   x"DA",   x"B1",   x"A4",   x"9B",   x"8E", 
  x"4D",   x"58",   x"67",   x"72",   x"19",   x"0C",   x"33",   x"26", 
  x"76",   x"63",   x"5C",   x"49",   x"22",   x"37",   x"08",   x"1D", 
  x"DE",   x"CB",   x"F4",   x"E1",   x"8A",   x"9F",   x"A0",   x"B5", 
  x"09",   x"1C",   x"23",   x"36",   x"5D",   x"48",   x"77",   x"62", 
  x"A1",   x"B4",   x"8B",   x"9E",   x"F5",   x"E0",   x"DF",   x"CA", 
  x"9A",   x"8F",   x"B0",   x"A5",   x"CE",   x"DB",   x"E4",   x"F1", 
  x"32",   x"27",   x"18",   x"0D",   x"66",   x"73",   x"4C",   x"59", 
  x"EC",   x"F9",   x"C6",   x"D3",   x"B8",   x"AD",   x"92",   x"87", 
  x"44",   x"51",   x"6E",   x"7B",   x"10",   x"05",   x"3A",   x"2F", 
  x"7F",   x"6A",   x"55",   x"40",   x"2B",   x"3E",   x"01",   x"14", 
  x"D7",   x"C2",   x"FD",   x"E8",   x"83",   x"96",   x"A9",   x"BC", 
  x"12",   x"07",   x"38",   x"2D",   x"46",   x"53",   x"6C",   x"79", 
  x"BA",   x"AF",   x"90",   x"85",   x"EE",   x"FB",   x"C4",   x"D1", 
  x"81",   x"94",   x"AB",   x"BE",   x"D5",   x"C0",   x"FF",   x"EA", 
  x"29",   x"3C",   x"03",   x"16",   x"7D",   x"68",   x"57",   x"42", 
  x"F7",   x"E2",   x"DD",   x"C8",   x"A3",   x"B6",   x"89",   x"9C", 
  x"5F",   x"4A",   x"75",   x"60",   x"0B",   x"1E",   x"21",   x"34", 
  x"64",   x"71",   x"4E",   x"5B",   x"30",   x"25",   x"1A",   x"0F", 
  x"CC",   x"D9",   x"E6",   x"F3",   x"98",   x"8D",   x"B2",   x"A7", 
  x"1B",   x"0E",   x"31",   x"24",   x"4F",   x"5A",   x"65",   x"70", 
  x"B3",   x"A6",   x"99",   x"8C",   x"E7",   x"F2",   x"CD",   x"D8", 
  x"88",   x"9D",   x"A2",   x"B7",   x"DC",   x"C9",   x"F6",   x"E3", 
  x"20",   x"35",   x"0A",   x"1F",   x"74",   x"61",   x"5E",   x"4B", 
  x"FE",   x"EB",   x"D4",   x"C1",   x"AA",   x"BF",   x"80",   x"95", 
  x"56",   x"43",   x"7C",   x"69",   x"02",   x"17",   x"28",   x"3D", 
  x"6D",   x"78",   x"47",   x"52",   x"39",   x"2C",   x"13",   x"06", 
  x"C5",   x"D0",   x"EF",   x"FA",   x"91",   x"84",   x"BB",   x"AE", 
  x"00",   x"16",   x"2C",   x"3A",   x"58",   x"4E",   x"74",   x"62", 
  x"B0",   x"A6",   x"9C",   x"8A",   x"E8",   x"FE",   x"C4",   x"D2", 
  x"A3",   x"B5",   x"8F",   x"99",   x"FB",   x"ED",   x"D7",   x"C1", 
  x"13",   x"05",   x"3F",   x"29",   x"4B",   x"5D",   x"67",   x"71", 
  x"85",   x"93",   x"A9",   x"BF",   x"DD",   x"CB",   x"F1",   x"E7", 
  x"35",   x"23",   x"19",   x"0F",   x"6D",   x"7B",   x"41",   x"57", 
  x"26",   x"30",   x"0A",   x"1C",   x"7E",   x"68",   x"52",   x"44", 
  x"96",   x"80",   x"BA",   x"AC",   x"CE",   x"D8",   x"E2",   x"F4", 
  x"C9",   x"DF",   x"E5",   x"F3",   x"91",   x"87",   x"BD",   x"AB", 
  x"79",   x"6F",   x"55",   x"43",   x"21",   x"37",   x"0D",   x"1B", 
  x"6A",   x"7C",   x"46",   x"50",   x"32",   x"24",   x"1E",   x"08", 
  x"DA",   x"CC",   x"F6",   x"E0",   x"82",   x"94",   x"AE",   x"B8", 
  x"4C",   x"5A",   x"60",   x"76",   x"14",   x"02",   x"38",   x"2E", 
  x"FC",   x"EA",   x"D0",   x"C6",   x"A4",   x"B2",   x"88",   x"9E", 
  x"EF",   x"F9",   x"C3",   x"D5",   x"B7",   x"A1",   x"9B",   x"8D", 
  x"5F",   x"49",   x"73",   x"65",   x"07",   x"11",   x"2B",   x"3D", 
  x"51",   x"47",   x"7D",   x"6B",   x"09",   x"1F",   x"25",   x"33", 
  x"E1",   x"F7",   x"CD",   x"DB",   x"B9",   x"AF",   x"95",   x"83", 
  x"F2",   x"E4",   x"DE",   x"C8",   x"AA",   x"BC",   x"86",   x"90", 
  x"42",   x"54",   x"6E",   x"78",   x"1A",   x"0C",   x"36",   x"20", 
  x"D4",   x"C2",   x"F8",   x"EE",   x"8C",   x"9A",   x"A0",   x"B6", 
  x"64",   x"72",   x"48",   x"5E",   x"3C",   x"2A",   x"10",   x"06", 
  x"77",   x"61",   x"5B",   x"4D",   x"2F",   x"39",   x"03",   x"15", 
  x"C7",   x"D1",   x"EB",   x"FD",   x"9F",   x"89",   x"B3",   x"A5", 
  x"98",   x"8E",   x"B4",   x"A2",   x"C0",   x"D6",   x"EC",   x"FA", 
  x"28",   x"3E",   x"04",   x"12",   x"70",   x"66",   x"5C",   x"4A", 
  x"3B",   x"2D",   x"17",   x"01",   x"63",   x"75",   x"4F",   x"59", 
  x"8B",   x"9D",   x"A7",   x"B1",   x"D3",   x"C5",   x"FF",   x"E9", 
  x"1D",   x"0B",   x"31",   x"27",   x"45",   x"53",   x"69",   x"7F", 
  x"AD",   x"BB",   x"81",   x"97",   x"F5",   x"E3",   x"D9",   x"CF", 
  x"BE",   x"A8",   x"92",   x"84",   x"E6",   x"F0",   x"CA",   x"DC", 
  x"0E",   x"18",   x"22",   x"34",   x"56",   x"40",   x"7A",   x"6C", 
  x"00",   x"17",   x"2E",   x"39",   x"5C",   x"4B",   x"72",   x"65", 
  x"B8",   x"AF",   x"96",   x"81",   x"E4",   x"F3",   x"CA",   x"DD", 
  x"B3",   x"A4",   x"9D",   x"8A",   x"EF",   x"F8",   x"C1",   x"D6", 
  x"0B",   x"1C",   x"25",   x"32",   x"57",   x"40",   x"79",   x"6E", 
  x"A5",   x"B2",   x"8B",   x"9C",   x"F9",   x"EE",   x"D7",   x"C0", 
  x"1D",   x"0A",   x"33",   x"24",   x"41",   x"56",   x"6F",   x"78", 
  x"16",   x"01",   x"38",   x"2F",   x"4A",   x"5D",   x"64",   x"73", 
  x"AE",   x"B9",   x"80",   x"97",   x"F2",   x"E5",   x"DC",   x"CB", 
  x"89",   x"9E",   x"A7",   x"B0",   x"D5",   x"C2",   x"FB",   x"EC", 
  x"31",   x"26",   x"1F",   x"08",   x"6D",   x"7A",   x"43",   x"54", 
  x"3A",   x"2D",   x"14",   x"03",   x"66",   x"71",   x"48",   x"5F", 
  x"82",   x"95",   x"AC",   x"BB",   x"DE",   x"C9",   x"F0",   x"E7", 
  x"2C",   x"3B",   x"02",   x"15",   x"70",   x"67",   x"5E",   x"49", 
  x"94",   x"83",   x"BA",   x"AD",   x"C8",   x"DF",   x"E6",   x"F1", 
  x"9F",   x"88",   x"B1",   x"A6",   x"C3",   x"D4",   x"ED",   x"FA", 
  x"27",   x"30",   x"09",   x"1E",   x"7B",   x"6C",   x"55",   x"42", 
  x"D1",   x"C6",   x"FF",   x"E8",   x"8D",   x"9A",   x"A3",   x"B4", 
  x"69",   x"7E",   x"47",   x"50",   x"35",   x"22",   x"1B",   x"0C", 
  x"62",   x"75",   x"4C",   x"5B",   x"3E",   x"29",   x"10",   x"07", 
  x"DA",   x"CD",   x"F4",   x"E3",   x"86",   x"91",   x"A8",   x"BF", 
  x"74",   x"63",   x"5A",   x"4D",   x"28",   x"3F",   x"06",   x"11", 
  x"CC",   x"DB",   x"E2",   x"F5",   x"90",   x"87",   x"BE",   x"A9", 
  x"C7",   x"D0",   x"E9",   x"FE",   x"9B",   x"8C",   x"B5",   x"A2", 
  x"7F",   x"68",   x"51",   x"46",   x"23",   x"34",   x"0D",   x"1A", 
  x"58",   x"4F",   x"76",   x"61",   x"04",   x"13",   x"2A",   x"3D", 
  x"E0",   x"F7",   x"CE",   x"D9",   x"BC",   x"AB",   x"92",   x"85", 
  x"EB",   x"FC",   x"C5",   x"D2",   x"B7",   x"A0",   x"99",   x"8E", 
  x"53",   x"44",   x"7D",   x"6A",   x"0F",   x"18",   x"21",   x"36", 
  x"FD",   x"EA",   x"D3",   x"C4",   x"A1",   x"B6",   x"8F",   x"98", 
  x"45",   x"52",   x"6B",   x"7C",   x"19",   x"0E",   x"37",   x"20", 
  x"4E",   x"59",   x"60",   x"77",   x"12",   x"05",   x"3C",   x"2B", 
  x"F6",   x"E1",   x"D8",   x"CF",   x"AA",   x"BD",   x"84",   x"93", 
  x"00",   x"18",   x"30",   x"28",   x"60",   x"78",   x"50",   x"48", 
  x"C0",   x"D8",   x"F0",   x"E8",   x"A0",   x"B8",   x"90",   x"88", 
  x"43",   x"5B",   x"73",   x"6B",   x"23",   x"3B",   x"13",   x"0B", 
  x"83",   x"9B",   x"B3",   x"AB",   x"E3",   x"FB",   x"D3",   x"CB", 
  x"86",   x"9E",   x"B6",   x"AE",   x"E6",   x"FE",   x"D6",   x"CE", 
  x"46",   x"5E",   x"76",   x"6E",   x"26",   x"3E",   x"16",   x"0E", 
  x"C5",   x"DD",   x"F5",   x"ED",   x"A5",   x"BD",   x"95",   x"8D", 
  x"05",   x"1D",   x"35",   x"2D",   x"65",   x"7D",   x"55",   x"4D", 
  x"CF",   x"D7",   x"FF",   x"E7",   x"AF",   x"B7",   x"9F",   x"87", 
  x"0F",   x"17",   x"3F",   x"27",   x"6F",   x"77",   x"5F",   x"47", 
  x"8C",   x"94",   x"BC",   x"A4",   x"EC",   x"F4",   x"DC",   x"C4", 
  x"4C",   x"54",   x"7C",   x"64",   x"2C",   x"34",   x"1C",   x"04", 
  x"49",   x"51",   x"79",   x"61",   x"29",   x"31",   x"19",   x"01", 
  x"89",   x"91",   x"B9",   x"A1",   x"E9",   x"F1",   x"D9",   x"C1", 
  x"0A",   x"12",   x"3A",   x"22",   x"6A",   x"72",   x"5A",   x"42", 
  x"CA",   x"D2",   x"FA",   x"E2",   x"AA",   x"B2",   x"9A",   x"82", 
  x"5D",   x"45",   x"6D",   x"75",   x"3D",   x"25",   x"0D",   x"15", 
  x"9D",   x"85",   x"AD",   x"B5",   x"FD",   x"E5",   x"CD",   x"D5", 
  x"1E",   x"06",   x"2E",   x"36",   x"7E",   x"66",   x"4E",   x"56", 
  x"DE",   x"C6",   x"EE",   x"F6",   x"BE",   x"A6",   x"8E",   x"96", 
  x"DB",   x"C3",   x"EB",   x"F3",   x"BB",   x"A3",   x"8B",   x"93", 
  x"1B",   x"03",   x"2B",   x"33",   x"7B",   x"63",   x"4B",   x"53", 
  x"98",   x"80",   x"A8",   x"B0",   x"F8",   x"E0",   x"C8",   x"D0", 
  x"58",   x"40",   x"68",   x"70",   x"38",   x"20",   x"08",   x"10", 
  x"92",   x"8A",   x"A2",   x"BA",   x"F2",   x"EA",   x"C2",   x"DA", 
  x"52",   x"4A",   x"62",   x"7A",   x"32",   x"2A",   x"02",   x"1A", 
  x"D1",   x"C9",   x"E1",   x"F9",   x"B1",   x"A9",   x"81",   x"99", 
  x"11",   x"09",   x"21",   x"39",   x"71",   x"69",   x"41",   x"59", 
  x"14",   x"0C",   x"24",   x"3C",   x"74",   x"6C",   x"44",   x"5C", 
  x"D4",   x"CC",   x"E4",   x"FC",   x"B4",   x"AC",   x"84",   x"9C", 
  x"57",   x"4F",   x"67",   x"7F",   x"37",   x"2F",   x"07",   x"1F", 
  x"97",   x"8F",   x"A7",   x"BF",   x"F7",   x"EF",   x"C7",   x"DF", 
  x"00",   x"19",   x"32",   x"2B",   x"64",   x"7D",   x"56",   x"4F", 
  x"C8",   x"D1",   x"FA",   x"E3",   x"AC",   x"B5",   x"9E",   x"87", 
  x"53",   x"4A",   x"61",   x"78",   x"37",   x"2E",   x"05",   x"1C", 
  x"9B",   x"82",   x"A9",   x"B0",   x"FF",   x"E6",   x"CD",   x"D4", 
  x"A6",   x"BF",   x"94",   x"8D",   x"C2",   x"DB",   x"F0",   x"E9", 
  x"6E",   x"77",   x"5C",   x"45",   x"0A",   x"13",   x"38",   x"21", 
  x"F5",   x"EC",   x"C7",   x"DE",   x"91",   x"88",   x"A3",   x"BA", 
  x"3D",   x"24",   x"0F",   x"16",   x"59",   x"40",   x"6B",   x"72", 
  x"8F",   x"96",   x"BD",   x"A4",   x"EB",   x"F2",   x"D9",   x"C0", 
  x"47",   x"5E",   x"75",   x"6C",   x"23",   x"3A",   x"11",   x"08", 
  x"DC",   x"C5",   x"EE",   x"F7",   x"B8",   x"A1",   x"8A",   x"93", 
  x"14",   x"0D",   x"26",   x"3F",   x"70",   x"69",   x"42",   x"5B", 
  x"29",   x"30",   x"1B",   x"02",   x"4D",   x"54",   x"7F",   x"66", 
  x"E1",   x"F8",   x"D3",   x"CA",   x"85",   x"9C",   x"B7",   x"AE", 
  x"7A",   x"63",   x"48",   x"51",   x"1E",   x"07",   x"2C",   x"35", 
  x"B2",   x"AB",   x"80",   x"99",   x"D6",   x"CF",   x"E4",   x"FD", 
  x"DD",   x"C4",   x"EF",   x"F6",   x"B9",   x"A0",   x"8B",   x"92", 
  x"15",   x"0C",   x"27",   x"3E",   x"71",   x"68",   x"43",   x"5A", 
  x"8E",   x"97",   x"BC",   x"A5",   x"EA",   x"F3",   x"D8",   x"C1", 
  x"46",   x"5F",   x"74",   x"6D",   x"22",   x"3B",   x"10",   x"09", 
  x"7B",   x"62",   x"49",   x"50",   x"1F",   x"06",   x"2D",   x"34", 
  x"B3",   x"AA",   x"81",   x"98",   x"D7",   x"CE",   x"E5",   x"FC", 
  x"28",   x"31",   x"1A",   x"03",   x"4C",   x"55",   x"7E",   x"67", 
  x"E0",   x"F9",   x"D2",   x"CB",   x"84",   x"9D",   x"B6",   x"AF", 
  x"52",   x"4B",   x"60",   x"79",   x"36",   x"2F",   x"04",   x"1D", 
  x"9A",   x"83",   x"A8",   x"B1",   x"FE",   x"E7",   x"CC",   x"D5", 
  x"01",   x"18",   x"33",   x"2A",   x"65",   x"7C",   x"57",   x"4E", 
  x"C9",   x"D0",   x"FB",   x"E2",   x"AD",   x"B4",   x"9F",   x"86", 
  x"F4",   x"ED",   x"C6",   x"DF",   x"90",   x"89",   x"A2",   x"BB", 
  x"3C",   x"25",   x"0E",   x"17",   x"58",   x"41",   x"6A",   x"73", 
  x"A7",   x"BE",   x"95",   x"8C",   x"C3",   x"DA",   x"F1",   x"E8", 
  x"6F",   x"76",   x"5D",   x"44",   x"0B",   x"12",   x"39",   x"20", 
  x"00",   x"1A",   x"34",   x"2E",   x"68",   x"72",   x"5C",   x"46", 
  x"D0",   x"CA",   x"E4",   x"FE",   x"B8",   x"A2",   x"8C",   x"96", 
  x"63",   x"79",   x"57",   x"4D",   x"0B",   x"11",   x"3F",   x"25", 
  x"B3",   x"A9",   x"87",   x"9D",   x"DB",   x"C1",   x"EF",   x"F5", 
  x"C6",   x"DC",   x"F2",   x"E8",   x"AE",   x"B4",   x"9A",   x"80", 
  x"16",   x"0C",   x"22",   x"38",   x"7E",   x"64",   x"4A",   x"50", 
  x"A5",   x"BF",   x"91",   x"8B",   x"CD",   x"D7",   x"F9",   x"E3", 
  x"75",   x"6F",   x"41",   x"5B",   x"1D",   x"07",   x"29",   x"33", 
  x"4F",   x"55",   x"7B",   x"61",   x"27",   x"3D",   x"13",   x"09", 
  x"9F",   x"85",   x"AB",   x"B1",   x"F7",   x"ED",   x"C3",   x"D9", 
  x"2C",   x"36",   x"18",   x"02",   x"44",   x"5E",   x"70",   x"6A", 
  x"FC",   x"E6",   x"C8",   x"D2",   x"94",   x"8E",   x"A0",   x"BA", 
  x"89",   x"93",   x"BD",   x"A7",   x"E1",   x"FB",   x"D5",   x"CF", 
  x"59",   x"43",   x"6D",   x"77",   x"31",   x"2B",   x"05",   x"1F", 
  x"EA",   x"F0",   x"DE",   x"C4",   x"82",   x"98",   x"B6",   x"AC", 
  x"3A",   x"20",   x"0E",   x"14",   x"52",   x"48",   x"66",   x"7C", 
  x"9E",   x"84",   x"AA",   x"B0",   x"F6",   x"EC",   x"C2",   x"D8", 
  x"4E",   x"54",   x"7A",   x"60",   x"26",   x"3C",   x"12",   x"08", 
  x"FD",   x"E7",   x"C9",   x"D3",   x"95",   x"8F",   x"A1",   x"BB", 
  x"2D",   x"37",   x"19",   x"03",   x"45",   x"5F",   x"71",   x"6B", 
  x"58",   x"42",   x"6C",   x"76",   x"30",   x"2A",   x"04",   x"1E", 
  x"88",   x"92",   x"BC",   x"A6",   x"E0",   x"FA",   x"D4",   x"CE", 
  x"3B",   x"21",   x"0F",   x"15",   x"53",   x"49",   x"67",   x"7D", 
  x"EB",   x"F1",   x"DF",   x"C5",   x"83",   x"99",   x"B7",   x"AD", 
  x"D1",   x"CB",   x"E5",   x"FF",   x"B9",   x"A3",   x"8D",   x"97", 
  x"01",   x"1B",   x"35",   x"2F",   x"69",   x"73",   x"5D",   x"47", 
  x"B2",   x"A8",   x"86",   x"9C",   x"DA",   x"C0",   x"EE",   x"F4", 
  x"62",   x"78",   x"56",   x"4C",   x"0A",   x"10",   x"3E",   x"24", 
  x"17",   x"0D",   x"23",   x"39",   x"7F",   x"65",   x"4B",   x"51", 
  x"C7",   x"DD",   x"F3",   x"E9",   x"AF",   x"B5",   x"9B",   x"81", 
  x"74",   x"6E",   x"40",   x"5A",   x"1C",   x"06",   x"28",   x"32", 
  x"A4",   x"BE",   x"90",   x"8A",   x"CC",   x"D6",   x"F8",   x"E2", 
  x"00",   x"1B",   x"36",   x"2D",   x"6C",   x"77",   x"5A",   x"41", 
  x"D8",   x"C3",   x"EE",   x"F5",   x"B4",   x"AF",   x"82",   x"99", 
  x"73",   x"68",   x"45",   x"5E",   x"1F",   x"04",   x"29",   x"32", 
  x"AB",   x"B0",   x"9D",   x"86",   x"C7",   x"DC",   x"F1",   x"EA", 
  x"E6",   x"FD",   x"D0",   x"CB",   x"8A",   x"91",   x"BC",   x"A7", 
  x"3E",   x"25",   x"08",   x"13",   x"52",   x"49",   x"64",   x"7F", 
  x"95",   x"8E",   x"A3",   x"B8",   x"F9",   x"E2",   x"CF",   x"D4", 
  x"4D",   x"56",   x"7B",   x"60",   x"21",   x"3A",   x"17",   x"0C", 
  x"0F",   x"14",   x"39",   x"22",   x"63",   x"78",   x"55",   x"4E", 
  x"D7",   x"CC",   x"E1",   x"FA",   x"BB",   x"A0",   x"8D",   x"96", 
  x"7C",   x"67",   x"4A",   x"51",   x"10",   x"0B",   x"26",   x"3D", 
  x"A4",   x"BF",   x"92",   x"89",   x"C8",   x"D3",   x"FE",   x"E5", 
  x"E9",   x"F2",   x"DF",   x"C4",   x"85",   x"9E",   x"B3",   x"A8", 
  x"31",   x"2A",   x"07",   x"1C",   x"5D",   x"46",   x"6B",   x"70", 
  x"9A",   x"81",   x"AC",   x"B7",   x"F6",   x"ED",   x"C0",   x"DB", 
  x"42",   x"59",   x"74",   x"6F",   x"2E",   x"35",   x"18",   x"03", 
  x"1E",   x"05",   x"28",   x"33",   x"72",   x"69",   x"44",   x"5F", 
  x"C6",   x"DD",   x"F0",   x"EB",   x"AA",   x"B1",   x"9C",   x"87", 
  x"6D",   x"76",   x"5B",   x"40",   x"01",   x"1A",   x"37",   x"2C", 
  x"B5",   x"AE",   x"83",   x"98",   x"D9",   x"C2",   x"EF",   x"F4", 
  x"F8",   x"E3",   x"CE",   x"D5",   x"94",   x"8F",   x"A2",   x"B9", 
  x"20",   x"3B",   x"16",   x"0D",   x"4C",   x"57",   x"7A",   x"61", 
  x"8B",   x"90",   x"BD",   x"A6",   x"E7",   x"FC",   x"D1",   x"CA", 
  x"53",   x"48",   x"65",   x"7E",   x"3F",   x"24",   x"09",   x"12", 
  x"11",   x"0A",   x"27",   x"3C",   x"7D",   x"66",   x"4B",   x"50", 
  x"C9",   x"D2",   x"FF",   x"E4",   x"A5",   x"BE",   x"93",   x"88", 
  x"62",   x"79",   x"54",   x"4F",   x"0E",   x"15",   x"38",   x"23", 
  x"BA",   x"A1",   x"8C",   x"97",   x"D6",   x"CD",   x"E0",   x"FB", 
  x"F7",   x"EC",   x"C1",   x"DA",   x"9B",   x"80",   x"AD",   x"B6", 
  x"2F",   x"34",   x"19",   x"02",   x"43",   x"58",   x"75",   x"6E", 
  x"84",   x"9F",   x"B2",   x"A9",   x"E8",   x"F3",   x"DE",   x"C5", 
  x"5C",   x"47",   x"6A",   x"71",   x"30",   x"2B",   x"06",   x"1D", 
  x"00",   x"1C",   x"38",   x"24",   x"70",   x"6C",   x"48",   x"54", 
  x"E0",   x"FC",   x"D8",   x"C4",   x"90",   x"8C",   x"A8",   x"B4", 
  x"03",   x"1F",   x"3B",   x"27",   x"73",   x"6F",   x"4B",   x"57", 
  x"E3",   x"FF",   x"DB",   x"C7",   x"93",   x"8F",   x"AB",   x"B7", 
  x"06",   x"1A",   x"3E",   x"22",   x"76",   x"6A",   x"4E",   x"52", 
  x"E6",   x"FA",   x"DE",   x"C2",   x"96",   x"8A",   x"AE",   x"B2", 
  x"05",   x"19",   x"3D",   x"21",   x"75",   x"69",   x"4D",   x"51", 
  x"E5",   x"F9",   x"DD",   x"C1",   x"95",   x"89",   x"AD",   x"B1", 
  x"0C",   x"10",   x"34",   x"28",   x"7C",   x"60",   x"44",   x"58", 
  x"EC",   x"F0",   x"D4",   x"C8",   x"9C",   x"80",   x"A4",   x"B8", 
  x"0F",   x"13",   x"37",   x"2B",   x"7F",   x"63",   x"47",   x"5B", 
  x"EF",   x"F3",   x"D7",   x"CB",   x"9F",   x"83",   x"A7",   x"BB", 
  x"0A",   x"16",   x"32",   x"2E",   x"7A",   x"66",   x"42",   x"5E", 
  x"EA",   x"F6",   x"D2",   x"CE",   x"9A",   x"86",   x"A2",   x"BE", 
  x"09",   x"15",   x"31",   x"2D",   x"79",   x"65",   x"41",   x"5D", 
  x"E9",   x"F5",   x"D1",   x"CD",   x"99",   x"85",   x"A1",   x"BD", 
  x"18",   x"04",   x"20",   x"3C",   x"68",   x"74",   x"50",   x"4C", 
  x"F8",   x"E4",   x"C0",   x"DC",   x"88",   x"94",   x"B0",   x"AC", 
  x"1B",   x"07",   x"23",   x"3F",   x"6B",   x"77",   x"53",   x"4F", 
  x"FB",   x"E7",   x"C3",   x"DF",   x"8B",   x"97",   x"B3",   x"AF", 
  x"1E",   x"02",   x"26",   x"3A",   x"6E",   x"72",   x"56",   x"4A", 
  x"FE",   x"E2",   x"C6",   x"DA",   x"8E",   x"92",   x"B6",   x"AA", 
  x"1D",   x"01",   x"25",   x"39",   x"6D",   x"71",   x"55",   x"49", 
  x"FD",   x"E1",   x"C5",   x"D9",   x"8D",   x"91",   x"B5",   x"A9", 
  x"14",   x"08",   x"2C",   x"30",   x"64",   x"78",   x"5C",   x"40", 
  x"F4",   x"E8",   x"CC",   x"D0",   x"84",   x"98",   x"BC",   x"A0", 
  x"17",   x"0B",   x"2F",   x"33",   x"67",   x"7B",   x"5F",   x"43", 
  x"F7",   x"EB",   x"CF",   x"D3",   x"87",   x"9B",   x"BF",   x"A3", 
  x"12",   x"0E",   x"2A",   x"36",   x"62",   x"7E",   x"5A",   x"46", 
  x"F2",   x"EE",   x"CA",   x"D6",   x"82",   x"9E",   x"BA",   x"A6", 
  x"11",   x"0D",   x"29",   x"35",   x"61",   x"7D",   x"59",   x"45", 
  x"F1",   x"ED",   x"C9",   x"D5",   x"81",   x"9D",   x"B9",   x"A5", 
  x"00",   x"1D",   x"3A",   x"27",   x"74",   x"69",   x"4E",   x"53", 
  x"E8",   x"F5",   x"D2",   x"CF",   x"9C",   x"81",   x"A6",   x"BB", 
  x"13",   x"0E",   x"29",   x"34",   x"67",   x"7A",   x"5D",   x"40", 
  x"FB",   x"E6",   x"C1",   x"DC",   x"8F",   x"92",   x"B5",   x"A8", 
  x"26",   x"3B",   x"1C",   x"01",   x"52",   x"4F",   x"68",   x"75", 
  x"CE",   x"D3",   x"F4",   x"E9",   x"BA",   x"A7",   x"80",   x"9D", 
  x"35",   x"28",   x"0F",   x"12",   x"41",   x"5C",   x"7B",   x"66", 
  x"DD",   x"C0",   x"E7",   x"FA",   x"A9",   x"B4",   x"93",   x"8E", 
  x"4C",   x"51",   x"76",   x"6B",   x"38",   x"25",   x"02",   x"1F", 
  x"A4",   x"B9",   x"9E",   x"83",   x"D0",   x"CD",   x"EA",   x"F7", 
  x"5F",   x"42",   x"65",   x"78",   x"2B",   x"36",   x"11",   x"0C", 
  x"B7",   x"AA",   x"8D",   x"90",   x"C3",   x"DE",   x"F9",   x"E4", 
  x"6A",   x"77",   x"50",   x"4D",   x"1E",   x"03",   x"24",   x"39", 
  x"82",   x"9F",   x"B8",   x"A5",   x"F6",   x"EB",   x"CC",   x"D1", 
  x"79",   x"64",   x"43",   x"5E",   x"0D",   x"10",   x"37",   x"2A", 
  x"91",   x"8C",   x"AB",   x"B6",   x"E5",   x"F8",   x"DF",   x"C2", 
  x"98",   x"85",   x"A2",   x"BF",   x"EC",   x"F1",   x"D6",   x"CB", 
  x"70",   x"6D",   x"4A",   x"57",   x"04",   x"19",   x"3E",   x"23", 
  x"8B",   x"96",   x"B1",   x"AC",   x"FF",   x"E2",   x"C5",   x"D8", 
  x"63",   x"7E",   x"59",   x"44",   x"17",   x"0A",   x"2D",   x"30", 
  x"BE",   x"A3",   x"84",   x"99",   x"CA",   x"D7",   x"F0",   x"ED", 
  x"56",   x"4B",   x"6C",   x"71",   x"22",   x"3F",   x"18",   x"05", 
  x"AD",   x"B0",   x"97",   x"8A",   x"D9",   x"C4",   x"E3",   x"FE", 
  x"45",   x"58",   x"7F",   x"62",   x"31",   x"2C",   x"0B",   x"16", 
  x"D4",   x"C9",   x"EE",   x"F3",   x"A0",   x"BD",   x"9A",   x"87", 
  x"3C",   x"21",   x"06",   x"1B",   x"48",   x"55",   x"72",   x"6F", 
  x"C7",   x"DA",   x"FD",   x"E0",   x"B3",   x"AE",   x"89",   x"94", 
  x"2F",   x"32",   x"15",   x"08",   x"5B",   x"46",   x"61",   x"7C", 
  x"F2",   x"EF",   x"C8",   x"D5",   x"86",   x"9B",   x"BC",   x"A1", 
  x"1A",   x"07",   x"20",   x"3D",   x"6E",   x"73",   x"54",   x"49", 
  x"E1",   x"FC",   x"DB",   x"C6",   x"95",   x"88",   x"AF",   x"B2", 
  x"09",   x"14",   x"33",   x"2E",   x"7D",   x"60",   x"47",   x"5A", 
  x"00",   x"1E",   x"3C",   x"22",   x"78",   x"66",   x"44",   x"5A", 
  x"F0",   x"EE",   x"CC",   x"D2",   x"88",   x"96",   x"B4",   x"AA", 
  x"23",   x"3D",   x"1F",   x"01",   x"5B",   x"45",   x"67",   x"79", 
  x"D3",   x"CD",   x"EF",   x"F1",   x"AB",   x"B5",   x"97",   x"89", 
  x"46",   x"58",   x"7A",   x"64",   x"3E",   x"20",   x"02",   x"1C", 
  x"B6",   x"A8",   x"8A",   x"94",   x"CE",   x"D0",   x"F2",   x"EC", 
  x"65",   x"7B",   x"59",   x"47",   x"1D",   x"03",   x"21",   x"3F", 
  x"95",   x"8B",   x"A9",   x"B7",   x"ED",   x"F3",   x"D1",   x"CF", 
  x"8C",   x"92",   x"B0",   x"AE",   x"F4",   x"EA",   x"C8",   x"D6", 
  x"7C",   x"62",   x"40",   x"5E",   x"04",   x"1A",   x"38",   x"26", 
  x"AF",   x"B1",   x"93",   x"8D",   x"D7",   x"C9",   x"EB",   x"F5", 
  x"5F",   x"41",   x"63",   x"7D",   x"27",   x"39",   x"1B",   x"05", 
  x"CA",   x"D4",   x"F6",   x"E8",   x"B2",   x"AC",   x"8E",   x"90", 
  x"3A",   x"24",   x"06",   x"18",   x"42",   x"5C",   x"7E",   x"60", 
  x"E9",   x"F7",   x"D5",   x"CB",   x"91",   x"8F",   x"AD",   x"B3", 
  x"19",   x"07",   x"25",   x"3B",   x"61",   x"7F",   x"5D",   x"43", 
  x"DB",   x"C5",   x"E7",   x"F9",   x"A3",   x"BD",   x"9F",   x"81", 
  x"2B",   x"35",   x"17",   x"09",   x"53",   x"4D",   x"6F",   x"71", 
  x"F8",   x"E6",   x"C4",   x"DA",   x"80",   x"9E",   x"BC",   x"A2", 
  x"08",   x"16",   x"34",   x"2A",   x"70",   x"6E",   x"4C",   x"52", 
  x"9D",   x"83",   x"A1",   x"BF",   x"E5",   x"FB",   x"D9",   x"C7", 
  x"6D",   x"73",   x"51",   x"4F",   x"15",   x"0B",   x"29",   x"37", 
  x"BE",   x"A0",   x"82",   x"9C",   x"C6",   x"D8",   x"FA",   x"E4", 
  x"4E",   x"50",   x"72",   x"6C",   x"36",   x"28",   x"0A",   x"14", 
  x"57",   x"49",   x"6B",   x"75",   x"2F",   x"31",   x"13",   x"0D", 
  x"A7",   x"B9",   x"9B",   x"85",   x"DF",   x"C1",   x"E3",   x"FD", 
  x"74",   x"6A",   x"48",   x"56",   x"0C",   x"12",   x"30",   x"2E", 
  x"84",   x"9A",   x"B8",   x"A6",   x"FC",   x"E2",   x"C0",   x"DE", 
  x"11",   x"0F",   x"2D",   x"33",   x"69",   x"77",   x"55",   x"4B", 
  x"E1",   x"FF",   x"DD",   x"C3",   x"99",   x"87",   x"A5",   x"BB", 
  x"32",   x"2C",   x"0E",   x"10",   x"4A",   x"54",   x"76",   x"68", 
  x"C2",   x"DC",   x"FE",   x"E0",   x"BA",   x"A4",   x"86",   x"98", 
  x"00",   x"1F",   x"3E",   x"21",   x"7C",   x"63",   x"42",   x"5D", 
  x"F8",   x"E7",   x"C6",   x"D9",   x"84",   x"9B",   x"BA",   x"A5", 
  x"33",   x"2C",   x"0D",   x"12",   x"4F",   x"50",   x"71",   x"6E", 
  x"CB",   x"D4",   x"F5",   x"EA",   x"B7",   x"A8",   x"89",   x"96", 
  x"66",   x"79",   x"58",   x"47",   x"1A",   x"05",   x"24",   x"3B", 
  x"9E",   x"81",   x"A0",   x"BF",   x"E2",   x"FD",   x"DC",   x"C3", 
  x"55",   x"4A",   x"6B",   x"74",   x"29",   x"36",   x"17",   x"08", 
  x"AD",   x"B2",   x"93",   x"8C",   x"D1",   x"CE",   x"EF",   x"F0", 
  x"CC",   x"D3",   x"F2",   x"ED",   x"B0",   x"AF",   x"8E",   x"91", 
  x"34",   x"2B",   x"0A",   x"15",   x"48",   x"57",   x"76",   x"69", 
  x"FF",   x"E0",   x"C1",   x"DE",   x"83",   x"9C",   x"BD",   x"A2", 
  x"07",   x"18",   x"39",   x"26",   x"7B",   x"64",   x"45",   x"5A", 
  x"AA",   x"B5",   x"94",   x"8B",   x"D6",   x"C9",   x"E8",   x"F7", 
  x"52",   x"4D",   x"6C",   x"73",   x"2E",   x"31",   x"10",   x"0F", 
  x"99",   x"86",   x"A7",   x"B8",   x"E5",   x"FA",   x"DB",   x"C4", 
  x"61",   x"7E",   x"5F",   x"40",   x"1D",   x"02",   x"23",   x"3C", 
  x"5B",   x"44",   x"65",   x"7A",   x"27",   x"38",   x"19",   x"06", 
  x"A3",   x"BC",   x"9D",   x"82",   x"DF",   x"C0",   x"E1",   x"FE", 
  x"68",   x"77",   x"56",   x"49",   x"14",   x"0B",   x"2A",   x"35", 
  x"90",   x"8F",   x"AE",   x"B1",   x"EC",   x"F3",   x"D2",   x"CD", 
  x"3D",   x"22",   x"03",   x"1C",   x"41",   x"5E",   x"7F",   x"60", 
  x"C5",   x"DA",   x"FB",   x"E4",   x"B9",   x"A6",   x"87",   x"98", 
  x"0E",   x"11",   x"30",   x"2F",   x"72",   x"6D",   x"4C",   x"53", 
  x"F6",   x"E9",   x"C8",   x"D7",   x"8A",   x"95",   x"B4",   x"AB", 
  x"97",   x"88",   x"A9",   x"B6",   x"EB",   x"F4",   x"D5",   x"CA", 
  x"6F",   x"70",   x"51",   x"4E",   x"13",   x"0C",   x"2D",   x"32", 
  x"A4",   x"BB",   x"9A",   x"85",   x"D8",   x"C7",   x"E6",   x"F9", 
  x"5C",   x"43",   x"62",   x"7D",   x"20",   x"3F",   x"1E",   x"01", 
  x"F1",   x"EE",   x"CF",   x"D0",   x"8D",   x"92",   x"B3",   x"AC", 
  x"09",   x"16",   x"37",   x"28",   x"75",   x"6A",   x"4B",   x"54", 
  x"C2",   x"DD",   x"FC",   x"E3",   x"BE",   x"A1",   x"80",   x"9F", 
  x"3A",   x"25",   x"04",   x"1B",   x"46",   x"59",   x"78",   x"67", 
  x"00",   x"20",   x"40",   x"60",   x"80",   x"A0",   x"C0",   x"E0", 
  x"C3",   x"E3",   x"83",   x"A3",   x"43",   x"63",   x"03",   x"23", 
  x"45",   x"65",   x"05",   x"25",   x"C5",   x"E5",   x"85",   x"A5", 
  x"86",   x"A6",   x"C6",   x"E6",   x"06",   x"26",   x"46",   x"66", 
  x"8A",   x"AA",   x"CA",   x"EA",   x"0A",   x"2A",   x"4A",   x"6A", 
  x"49",   x"69",   x"09",   x"29",   x"C9",   x"E9",   x"89",   x"A9", 
  x"CF",   x"EF",   x"8F",   x"AF",   x"4F",   x"6F",   x"0F",   x"2F", 
  x"0C",   x"2C",   x"4C",   x"6C",   x"8C",   x"AC",   x"CC",   x"EC", 
  x"D7",   x"F7",   x"97",   x"B7",   x"57",   x"77",   x"17",   x"37", 
  x"14",   x"34",   x"54",   x"74",   x"94",   x"B4",   x"D4",   x"F4", 
  x"92",   x"B2",   x"D2",   x"F2",   x"12",   x"32",   x"52",   x"72", 
  x"51",   x"71",   x"11",   x"31",   x"D1",   x"F1",   x"91",   x"B1", 
  x"5D",   x"7D",   x"1D",   x"3D",   x"DD",   x"FD",   x"9D",   x"BD", 
  x"9E",   x"BE",   x"DE",   x"FE",   x"1E",   x"3E",   x"5E",   x"7E", 
  x"18",   x"38",   x"58",   x"78",   x"98",   x"B8",   x"D8",   x"F8", 
  x"DB",   x"FB",   x"9B",   x"BB",   x"5B",   x"7B",   x"1B",   x"3B", 
  x"6D",   x"4D",   x"2D",   x"0D",   x"ED",   x"CD",   x"AD",   x"8D", 
  x"AE",   x"8E",   x"EE",   x"CE",   x"2E",   x"0E",   x"6E",   x"4E", 
  x"28",   x"08",   x"68",   x"48",   x"A8",   x"88",   x"E8",   x"C8", 
  x"EB",   x"CB",   x"AB",   x"8B",   x"6B",   x"4B",   x"2B",   x"0B", 
  x"E7",   x"C7",   x"A7",   x"87",   x"67",   x"47",   x"27",   x"07", 
  x"24",   x"04",   x"64",   x"44",   x"A4",   x"84",   x"E4",   x"C4", 
  x"A2",   x"82",   x"E2",   x"C2",   x"22",   x"02",   x"62",   x"42", 
  x"61",   x"41",   x"21",   x"01",   x"E1",   x"C1",   x"A1",   x"81", 
  x"BA",   x"9A",   x"FA",   x"DA",   x"3A",   x"1A",   x"7A",   x"5A", 
  x"79",   x"59",   x"39",   x"19",   x"F9",   x"D9",   x"B9",   x"99", 
  x"FF",   x"DF",   x"BF",   x"9F",   x"7F",   x"5F",   x"3F",   x"1F", 
  x"3C",   x"1C",   x"7C",   x"5C",   x"BC",   x"9C",   x"FC",   x"DC", 
  x"30",   x"10",   x"70",   x"50",   x"B0",   x"90",   x"F0",   x"D0", 
  x"F3",   x"D3",   x"B3",   x"93",   x"73",   x"53",   x"33",   x"13", 
  x"75",   x"55",   x"35",   x"15",   x"F5",   x"D5",   x"B5",   x"95", 
  x"B6",   x"96",   x"F6",   x"D6",   x"36",   x"16",   x"76",   x"56", 
  x"00",   x"21",   x"42",   x"63",   x"84",   x"A5",   x"C6",   x"E7", 
  x"CB",   x"EA",   x"89",   x"A8",   x"4F",   x"6E",   x"0D",   x"2C", 
  x"55",   x"74",   x"17",   x"36",   x"D1",   x"F0",   x"93",   x"B2", 
  x"9E",   x"BF",   x"DC",   x"FD",   x"1A",   x"3B",   x"58",   x"79", 
  x"AA",   x"8B",   x"E8",   x"C9",   x"2E",   x"0F",   x"6C",   x"4D", 
  x"61",   x"40",   x"23",   x"02",   x"E5",   x"C4",   x"A7",   x"86", 
  x"FF",   x"DE",   x"BD",   x"9C",   x"7B",   x"5A",   x"39",   x"18", 
  x"34",   x"15",   x"76",   x"57",   x"B0",   x"91",   x"F2",   x"D3", 
  x"97",   x"B6",   x"D5",   x"F4",   x"13",   x"32",   x"51",   x"70", 
  x"5C",   x"7D",   x"1E",   x"3F",   x"D8",   x"F9",   x"9A",   x"BB", 
  x"C2",   x"E3",   x"80",   x"A1",   x"46",   x"67",   x"04",   x"25", 
  x"09",   x"28",   x"4B",   x"6A",   x"8D",   x"AC",   x"CF",   x"EE", 
  x"3D",   x"1C",   x"7F",   x"5E",   x"B9",   x"98",   x"FB",   x"DA", 
  x"F6",   x"D7",   x"B4",   x"95",   x"72",   x"53",   x"30",   x"11", 
  x"68",   x"49",   x"2A",   x"0B",   x"EC",   x"CD",   x"AE",   x"8F", 
  x"A3",   x"82",   x"E1",   x"C0",   x"27",   x"06",   x"65",   x"44", 
  x"ED",   x"CC",   x"AF",   x"8E",   x"69",   x"48",   x"2B",   x"0A", 
  x"26",   x"07",   x"64",   x"45",   x"A2",   x"83",   x"E0",   x"C1", 
  x"B8",   x"99",   x"FA",   x"DB",   x"3C",   x"1D",   x"7E",   x"5F", 
  x"73",   x"52",   x"31",   x"10",   x"F7",   x"D6",   x"B5",   x"94", 
  x"47",   x"66",   x"05",   x"24",   x"C3",   x"E2",   x"81",   x"A0", 
  x"8C",   x"AD",   x"CE",   x"EF",   x"08",   x"29",   x"4A",   x"6B", 
  x"12",   x"33",   x"50",   x"71",   x"96",   x"B7",   x"D4",   x"F5", 
  x"D9",   x"F8",   x"9B",   x"BA",   x"5D",   x"7C",   x"1F",   x"3E", 
  x"7A",   x"5B",   x"38",   x"19",   x"FE",   x"DF",   x"BC",   x"9D", 
  x"B1",   x"90",   x"F3",   x"D2",   x"35",   x"14",   x"77",   x"56", 
  x"2F",   x"0E",   x"6D",   x"4C",   x"AB",   x"8A",   x"E9",   x"C8", 
  x"E4",   x"C5",   x"A6",   x"87",   x"60",   x"41",   x"22",   x"03", 
  x"D0",   x"F1",   x"92",   x"B3",   x"54",   x"75",   x"16",   x"37", 
  x"1B",   x"3A",   x"59",   x"78",   x"9F",   x"BE",   x"DD",   x"FC", 
  x"85",   x"A4",   x"C7",   x"E6",   x"01",   x"20",   x"43",   x"62", 
  x"4E",   x"6F",   x"0C",   x"2D",   x"CA",   x"EB",   x"88",   x"A9", 
  x"00",   x"22",   x"44",   x"66",   x"88",   x"AA",   x"CC",   x"EE", 
  x"D3",   x"F1",   x"97",   x"B5",   x"5B",   x"79",   x"1F",   x"3D", 
  x"65",   x"47",   x"21",   x"03",   x"ED",   x"CF",   x"A9",   x"8B", 
  x"B6",   x"94",   x"F2",   x"D0",   x"3E",   x"1C",   x"7A",   x"58", 
  x"CA",   x"E8",   x"8E",   x"AC",   x"42",   x"60",   x"06",   x"24", 
  x"19",   x"3B",   x"5D",   x"7F",   x"91",   x"B3",   x"D5",   x"F7", 
  x"AF",   x"8D",   x"EB",   x"C9",   x"27",   x"05",   x"63",   x"41", 
  x"7C",   x"5E",   x"38",   x"1A",   x"F4",   x"D6",   x"B0",   x"92", 
  x"57",   x"75",   x"13",   x"31",   x"DF",   x"FD",   x"9B",   x"B9", 
  x"84",   x"A6",   x"C0",   x"E2",   x"0C",   x"2E",   x"48",   x"6A", 
  x"32",   x"10",   x"76",   x"54",   x"BA",   x"98",   x"FE",   x"DC", 
  x"E1",   x"C3",   x"A5",   x"87",   x"69",   x"4B",   x"2D",   x"0F", 
  x"9D",   x"BF",   x"D9",   x"FB",   x"15",   x"37",   x"51",   x"73", 
  x"4E",   x"6C",   x"0A",   x"28",   x"C6",   x"E4",   x"82",   x"A0", 
  x"F8",   x"DA",   x"BC",   x"9E",   x"70",   x"52",   x"34",   x"16", 
  x"2B",   x"09",   x"6F",   x"4D",   x"A3",   x"81",   x"E7",   x"C5", 
  x"AE",   x"8C",   x"EA",   x"C8",   x"26",   x"04",   x"62",   x"40", 
  x"7D",   x"5F",   x"39",   x"1B",   x"F5",   x"D7",   x"B1",   x"93", 
  x"CB",   x"E9",   x"8F",   x"AD",   x"43",   x"61",   x"07",   x"25", 
  x"18",   x"3A",   x"5C",   x"7E",   x"90",   x"B2",   x"D4",   x"F6", 
  x"64",   x"46",   x"20",   x"02",   x"EC",   x"CE",   x"A8",   x"8A", 
  x"B7",   x"95",   x"F3",   x"D1",   x"3F",   x"1D",   x"7B",   x"59", 
  x"01",   x"23",   x"45",   x"67",   x"89",   x"AB",   x"CD",   x"EF", 
  x"D2",   x"F0",   x"96",   x"B4",   x"5A",   x"78",   x"1E",   x"3C", 
  x"F9",   x"DB",   x"BD",   x"9F",   x"71",   x"53",   x"35",   x"17", 
  x"2A",   x"08",   x"6E",   x"4C",   x"A2",   x"80",   x"E6",   x"C4", 
  x"9C",   x"BE",   x"D8",   x"FA",   x"14",   x"36",   x"50",   x"72", 
  x"4F",   x"6D",   x"0B",   x"29",   x"C7",   x"E5",   x"83",   x"A1", 
  x"33",   x"11",   x"77",   x"55",   x"BB",   x"99",   x"FF",   x"DD", 
  x"E0",   x"C2",   x"A4",   x"86",   x"68",   x"4A",   x"2C",   x"0E", 
  x"56",   x"74",   x"12",   x"30",   x"DE",   x"FC",   x"9A",   x"B8", 
  x"85",   x"A7",   x"C1",   x"E3",   x"0D",   x"2F",   x"49",   x"6B", 
  x"00",   x"23",   x"46",   x"65",   x"8C",   x"AF",   x"CA",   x"E9", 
  x"DB",   x"F8",   x"9D",   x"BE",   x"57",   x"74",   x"11",   x"32", 
  x"75",   x"56",   x"33",   x"10",   x"F9",   x"DA",   x"BF",   x"9C", 
  x"AE",   x"8D",   x"E8",   x"CB",   x"22",   x"01",   x"64",   x"47", 
  x"EA",   x"C9",   x"AC",   x"8F",   x"66",   x"45",   x"20",   x"03", 
  x"31",   x"12",   x"77",   x"54",   x"BD",   x"9E",   x"FB",   x"D8", 
  x"9F",   x"BC",   x"D9",   x"FA",   x"13",   x"30",   x"55",   x"76", 
  x"44",   x"67",   x"02",   x"21",   x"C8",   x"EB",   x"8E",   x"AD", 
  x"17",   x"34",   x"51",   x"72",   x"9B",   x"B8",   x"DD",   x"FE", 
  x"CC",   x"EF",   x"8A",   x"A9",   x"40",   x"63",   x"06",   x"25", 
  x"62",   x"41",   x"24",   x"07",   x"EE",   x"CD",   x"A8",   x"8B", 
  x"B9",   x"9A",   x"FF",   x"DC",   x"35",   x"16",   x"73",   x"50", 
  x"FD",   x"DE",   x"BB",   x"98",   x"71",   x"52",   x"37",   x"14", 
  x"26",   x"05",   x"60",   x"43",   x"AA",   x"89",   x"EC",   x"CF", 
  x"88",   x"AB",   x"CE",   x"ED",   x"04",   x"27",   x"42",   x"61", 
  x"53",   x"70",   x"15",   x"36",   x"DF",   x"FC",   x"99",   x"BA", 
  x"2E",   x"0D",   x"68",   x"4B",   x"A2",   x"81",   x"E4",   x"C7", 
  x"F5",   x"D6",   x"B3",   x"90",   x"79",   x"5A",   x"3F",   x"1C", 
  x"5B",   x"78",   x"1D",   x"3E",   x"D7",   x"F4",   x"91",   x"B2", 
  x"80",   x"A3",   x"C6",   x"E5",   x"0C",   x"2F",   x"4A",   x"69", 
  x"C4",   x"E7",   x"82",   x"A1",   x"48",   x"6B",   x"0E",   x"2D", 
  x"1F",   x"3C",   x"59",   x"7A",   x"93",   x"B0",   x"D5",   x"F6", 
  x"B1",   x"92",   x"F7",   x"D4",   x"3D",   x"1E",   x"7B",   x"58", 
  x"6A",   x"49",   x"2C",   x"0F",   x"E6",   x"C5",   x"A0",   x"83", 
  x"39",   x"1A",   x"7F",   x"5C",   x"B5",   x"96",   x"F3",   x"D0", 
  x"E2",   x"C1",   x"A4",   x"87",   x"6E",   x"4D",   x"28",   x"0B", 
  x"4C",   x"6F",   x"0A",   x"29",   x"C0",   x"E3",   x"86",   x"A5", 
  x"97",   x"B4",   x"D1",   x"F2",   x"1B",   x"38",   x"5D",   x"7E", 
  x"D3",   x"F0",   x"95",   x"B6",   x"5F",   x"7C",   x"19",   x"3A", 
  x"08",   x"2B",   x"4E",   x"6D",   x"84",   x"A7",   x"C2",   x"E1", 
  x"A6",   x"85",   x"E0",   x"C3",   x"2A",   x"09",   x"6C",   x"4F", 
  x"7D",   x"5E",   x"3B",   x"18",   x"F1",   x"D2",   x"B7",   x"94", 
  x"00",   x"24",   x"48",   x"6C",   x"90",   x"B4",   x"D8",   x"FC", 
  x"E3",   x"C7",   x"AB",   x"8F",   x"73",   x"57",   x"3B",   x"1F", 
  x"05",   x"21",   x"4D",   x"69",   x"95",   x"B1",   x"DD",   x"F9", 
  x"E6",   x"C2",   x"AE",   x"8A",   x"76",   x"52",   x"3E",   x"1A", 
  x"0A",   x"2E",   x"42",   x"66",   x"9A",   x"BE",   x"D2",   x"F6", 
  x"E9",   x"CD",   x"A1",   x"85",   x"79",   x"5D",   x"31",   x"15", 
  x"0F",   x"2B",   x"47",   x"63",   x"9F",   x"BB",   x"D7",   x"F3", 
  x"EC",   x"C8",   x"A4",   x"80",   x"7C",   x"58",   x"34",   x"10", 
  x"14",   x"30",   x"5C",   x"78",   x"84",   x"A0",   x"CC",   x"E8", 
  x"F7",   x"D3",   x"BF",   x"9B",   x"67",   x"43",   x"2F",   x"0B", 
  x"11",   x"35",   x"59",   x"7D",   x"81",   x"A5",   x"C9",   x"ED", 
  x"F2",   x"D6",   x"BA",   x"9E",   x"62",   x"46",   x"2A",   x"0E", 
  x"1E",   x"3A",   x"56",   x"72",   x"8E",   x"AA",   x"C6",   x"E2", 
  x"FD",   x"D9",   x"B5",   x"91",   x"6D",   x"49",   x"25",   x"01", 
  x"1B",   x"3F",   x"53",   x"77",   x"8B",   x"AF",   x"C3",   x"E7", 
  x"F8",   x"DC",   x"B0",   x"94",   x"68",   x"4C",   x"20",   x"04", 
  x"28",   x"0C",   x"60",   x"44",   x"B8",   x"9C",   x"F0",   x"D4", 
  x"CB",   x"EF",   x"83",   x"A7",   x"5B",   x"7F",   x"13",   x"37", 
  x"2D",   x"09",   x"65",   x"41",   x"BD",   x"99",   x"F5",   x"D1", 
  x"CE",   x"EA",   x"86",   x"A2",   x"5E",   x"7A",   x"16",   x"32", 
  x"22",   x"06",   x"6A",   x"4E",   x"B2",   x"96",   x"FA",   x"DE", 
  x"C1",   x"E5",   x"89",   x"AD",   x"51",   x"75",   x"19",   x"3D", 
  x"27",   x"03",   x"6F",   x"4B",   x"B7",   x"93",   x"FF",   x"DB", 
  x"C4",   x"E0",   x"8C",   x"A8",   x"54",   x"70",   x"1C",   x"38", 
  x"3C",   x"18",   x"74",   x"50",   x"AC",   x"88",   x"E4",   x"C0", 
  x"DF",   x"FB",   x"97",   x"B3",   x"4F",   x"6B",   x"07",   x"23", 
  x"39",   x"1D",   x"71",   x"55",   x"A9",   x"8D",   x"E1",   x"C5", 
  x"DA",   x"FE",   x"92",   x"B6",   x"4A",   x"6E",   x"02",   x"26", 
  x"36",   x"12",   x"7E",   x"5A",   x"A6",   x"82",   x"EE",   x"CA", 
  x"D5",   x"F1",   x"9D",   x"B9",   x"45",   x"61",   x"0D",   x"29", 
  x"33",   x"17",   x"7B",   x"5F",   x"A3",   x"87",   x"EB",   x"CF", 
  x"D0",   x"F4",   x"98",   x"BC",   x"40",   x"64",   x"08",   x"2C", 
  x"00",   x"25",   x"4A",   x"6F",   x"94",   x"B1",   x"DE",   x"FB", 
  x"EB",   x"CE",   x"A1",   x"84",   x"7F",   x"5A",   x"35",   x"10", 
  x"15",   x"30",   x"5F",   x"7A",   x"81",   x"A4",   x"CB",   x"EE", 
  x"FE",   x"DB",   x"B4",   x"91",   x"6A",   x"4F",   x"20",   x"05", 
  x"2A",   x"0F",   x"60",   x"45",   x"BE",   x"9B",   x"F4",   x"D1", 
  x"C1",   x"E4",   x"8B",   x"AE",   x"55",   x"70",   x"1F",   x"3A", 
  x"3F",   x"1A",   x"75",   x"50",   x"AB",   x"8E",   x"E1",   x"C4", 
  x"D4",   x"F1",   x"9E",   x"BB",   x"40",   x"65",   x"0A",   x"2F", 
  x"54",   x"71",   x"1E",   x"3B",   x"C0",   x"E5",   x"8A",   x"AF", 
  x"BF",   x"9A",   x"F5",   x"D0",   x"2B",   x"0E",   x"61",   x"44", 
  x"41",   x"64",   x"0B",   x"2E",   x"D5",   x"F0",   x"9F",   x"BA", 
  x"AA",   x"8F",   x"E0",   x"C5",   x"3E",   x"1B",   x"74",   x"51", 
  x"7E",   x"5B",   x"34",   x"11",   x"EA",   x"CF",   x"A0",   x"85", 
  x"95",   x"B0",   x"DF",   x"FA",   x"01",   x"24",   x"4B",   x"6E", 
  x"6B",   x"4E",   x"21",   x"04",   x"FF",   x"DA",   x"B5",   x"90", 
  x"80",   x"A5",   x"CA",   x"EF",   x"14",   x"31",   x"5E",   x"7B", 
  x"A8",   x"8D",   x"E2",   x"C7",   x"3C",   x"19",   x"76",   x"53", 
  x"43",   x"66",   x"09",   x"2C",   x"D7",   x"F2",   x"9D",   x"B8", 
  x"BD",   x"98",   x"F7",   x"D2",   x"29",   x"0C",   x"63",   x"46", 
  x"56",   x"73",   x"1C",   x"39",   x"C2",   x"E7",   x"88",   x"AD", 
  x"82",   x"A7",   x"C8",   x"ED",   x"16",   x"33",   x"5C",   x"79", 
  x"69",   x"4C",   x"23",   x"06",   x"FD",   x"D8",   x"B7",   x"92", 
  x"97",   x"B2",   x"DD",   x"F8",   x"03",   x"26",   x"49",   x"6C", 
  x"7C",   x"59",   x"36",   x"13",   x"E8",   x"CD",   x"A2",   x"87", 
  x"FC",   x"D9",   x"B6",   x"93",   x"68",   x"4D",   x"22",   x"07", 
  x"17",   x"32",   x"5D",   x"78",   x"83",   x"A6",   x"C9",   x"EC", 
  x"E9",   x"CC",   x"A3",   x"86",   x"7D",   x"58",   x"37",   x"12", 
  x"02",   x"27",   x"48",   x"6D",   x"96",   x"B3",   x"DC",   x"F9", 
  x"D6",   x"F3",   x"9C",   x"B9",   x"42",   x"67",   x"08",   x"2D", 
  x"3D",   x"18",   x"77",   x"52",   x"A9",   x"8C",   x"E3",   x"C6", 
  x"C3",   x"E6",   x"89",   x"AC",   x"57",   x"72",   x"1D",   x"38", 
  x"28",   x"0D",   x"62",   x"47",   x"BC",   x"99",   x"F6",   x"D3", 
  x"00",   x"26",   x"4C",   x"6A",   x"98",   x"BE",   x"D4",   x"F2", 
  x"F3",   x"D5",   x"BF",   x"99",   x"6B",   x"4D",   x"27",   x"01", 
  x"25",   x"03",   x"69",   x"4F",   x"BD",   x"9B",   x"F1",   x"D7", 
  x"D6",   x"F0",   x"9A",   x"BC",   x"4E",   x"68",   x"02",   x"24", 
  x"4A",   x"6C",   x"06",   x"20",   x"D2",   x"F4",   x"9E",   x"B8", 
  x"B9",   x"9F",   x"F5",   x"D3",   x"21",   x"07",   x"6D",   x"4B", 
  x"6F",   x"49",   x"23",   x"05",   x"F7",   x"D1",   x"BB",   x"9D", 
  x"9C",   x"BA",   x"D0",   x"F6",   x"04",   x"22",   x"48",   x"6E", 
  x"94",   x"B2",   x"D8",   x"FE",   x"0C",   x"2A",   x"40",   x"66", 
  x"67",   x"41",   x"2B",   x"0D",   x"FF",   x"D9",   x"B3",   x"95", 
  x"B1",   x"97",   x"FD",   x"DB",   x"29",   x"0F",   x"65",   x"43", 
  x"42",   x"64",   x"0E",   x"28",   x"DA",   x"FC",   x"96",   x"B0", 
  x"DE",   x"F8",   x"92",   x"B4",   x"46",   x"60",   x"0A",   x"2C", 
  x"2D",   x"0B",   x"61",   x"47",   x"B5",   x"93",   x"F9",   x"DF", 
  x"FB",   x"DD",   x"B7",   x"91",   x"63",   x"45",   x"2F",   x"09", 
  x"08",   x"2E",   x"44",   x"62",   x"90",   x"B6",   x"DC",   x"FA", 
  x"EB",   x"CD",   x"A7",   x"81",   x"73",   x"55",   x"3F",   x"19", 
  x"18",   x"3E",   x"54",   x"72",   x"80",   x"A6",   x"CC",   x"EA", 
  x"CE",   x"E8",   x"82",   x"A4",   x"56",   x"70",   x"1A",   x"3C", 
  x"3D",   x"1B",   x"71",   x"57",   x"A5",   x"83",   x"E9",   x"CF", 
  x"A1",   x"87",   x"ED",   x"CB",   x"39",   x"1F",   x"75",   x"53", 
  x"52",   x"74",   x"1E",   x"38",   x"CA",   x"EC",   x"86",   x"A0", 
  x"84",   x"A2",   x"C8",   x"EE",   x"1C",   x"3A",   x"50",   x"76", 
  x"77",   x"51",   x"3B",   x"1D",   x"EF",   x"C9",   x"A3",   x"85", 
  x"7F",   x"59",   x"33",   x"15",   x"E7",   x"C1",   x"AB",   x"8D", 
  x"8C",   x"AA",   x"C0",   x"E6",   x"14",   x"32",   x"58",   x"7E", 
  x"5A",   x"7C",   x"16",   x"30",   x"C2",   x"E4",   x"8E",   x"A8", 
  x"A9",   x"8F",   x"E5",   x"C3",   x"31",   x"17",   x"7D",   x"5B", 
  x"35",   x"13",   x"79",   x"5F",   x"AD",   x"8B",   x"E1",   x"C7", 
  x"C6",   x"E0",   x"8A",   x"AC",   x"5E",   x"78",   x"12",   x"34", 
  x"10",   x"36",   x"5C",   x"7A",   x"88",   x"AE",   x"C4",   x"E2", 
  x"E3",   x"C5",   x"AF",   x"89",   x"7B",   x"5D",   x"37",   x"11", 
  x"00",   x"27",   x"4E",   x"69",   x"9C",   x"BB",   x"D2",   x"F5", 
  x"FB",   x"DC",   x"B5",   x"92",   x"67",   x"40",   x"29",   x"0E", 
  x"35",   x"12",   x"7B",   x"5C",   x"A9",   x"8E",   x"E7",   x"C0", 
  x"CE",   x"E9",   x"80",   x"A7",   x"52",   x"75",   x"1C",   x"3B", 
  x"6A",   x"4D",   x"24",   x"03",   x"F6",   x"D1",   x"B8",   x"9F", 
  x"91",   x"B6",   x"DF",   x"F8",   x"0D",   x"2A",   x"43",   x"64", 
  x"5F",   x"78",   x"11",   x"36",   x"C3",   x"E4",   x"8D",   x"AA", 
  x"A4",   x"83",   x"EA",   x"CD",   x"38",   x"1F",   x"76",   x"51", 
  x"D4",   x"F3",   x"9A",   x"BD",   x"48",   x"6F",   x"06",   x"21", 
  x"2F",   x"08",   x"61",   x"46",   x"B3",   x"94",   x"FD",   x"DA", 
  x"E1",   x"C6",   x"AF",   x"88",   x"7D",   x"5A",   x"33",   x"14", 
  x"1A",   x"3D",   x"54",   x"73",   x"86",   x"A1",   x"C8",   x"EF", 
  x"BE",   x"99",   x"F0",   x"D7",   x"22",   x"05",   x"6C",   x"4B", 
  x"45",   x"62",   x"0B",   x"2C",   x"D9",   x"FE",   x"97",   x"B0", 
  x"8B",   x"AC",   x"C5",   x"E2",   x"17",   x"30",   x"59",   x"7E", 
  x"70",   x"57",   x"3E",   x"19",   x"EC",   x"CB",   x"A2",   x"85", 
  x"6B",   x"4C",   x"25",   x"02",   x"F7",   x"D0",   x"B9",   x"9E", 
  x"90",   x"B7",   x"DE",   x"F9",   x"0C",   x"2B",   x"42",   x"65", 
  x"5E",   x"79",   x"10",   x"37",   x"C2",   x"E5",   x"8C",   x"AB", 
  x"A5",   x"82",   x"EB",   x"CC",   x"39",   x"1E",   x"77",   x"50", 
  x"01",   x"26",   x"4F",   x"68",   x"9D",   x"BA",   x"D3",   x"F4", 
  x"FA",   x"DD",   x"B4",   x"93",   x"66",   x"41",   x"28",   x"0F", 
  x"34",   x"13",   x"7A",   x"5D",   x"A8",   x"8F",   x"E6",   x"C1", 
  x"CF",   x"E8",   x"81",   x"A6",   x"53",   x"74",   x"1D",   x"3A", 
  x"BF",   x"98",   x"F1",   x"D6",   x"23",   x"04",   x"6D",   x"4A", 
  x"44",   x"63",   x"0A",   x"2D",   x"D8",   x"FF",   x"96",   x"B1", 
  x"8A",   x"AD",   x"C4",   x"E3",   x"16",   x"31",   x"58",   x"7F", 
  x"71",   x"56",   x"3F",   x"18",   x"ED",   x"CA",   x"A3",   x"84", 
  x"D5",   x"F2",   x"9B",   x"BC",   x"49",   x"6E",   x"07",   x"20", 
  x"2E",   x"09",   x"60",   x"47",   x"B2",   x"95",   x"FC",   x"DB", 
  x"E0",   x"C7",   x"AE",   x"89",   x"7C",   x"5B",   x"32",   x"15", 
  x"1B",   x"3C",   x"55",   x"72",   x"87",   x"A0",   x"C9",   x"EE", 
  x"00",   x"28",   x"50",   x"78",   x"A0",   x"88",   x"F0",   x"D8", 
  x"83",   x"AB",   x"D3",   x"FB",   x"23",   x"0B",   x"73",   x"5B", 
  x"C5",   x"ED",   x"95",   x"BD",   x"65",   x"4D",   x"35",   x"1D", 
  x"46",   x"6E",   x"16",   x"3E",   x"E6",   x"CE",   x"B6",   x"9E", 
  x"49",   x"61",   x"19",   x"31",   x"E9",   x"C1",   x"B9",   x"91", 
  x"CA",   x"E2",   x"9A",   x"B2",   x"6A",   x"42",   x"3A",   x"12", 
  x"8C",   x"A4",   x"DC",   x"F4",   x"2C",   x"04",   x"7C",   x"54", 
  x"0F",   x"27",   x"5F",   x"77",   x"AF",   x"87",   x"FF",   x"D7", 
  x"92",   x"BA",   x"C2",   x"EA",   x"32",   x"1A",   x"62",   x"4A", 
  x"11",   x"39",   x"41",   x"69",   x"B1",   x"99",   x"E1",   x"C9", 
  x"57",   x"7F",   x"07",   x"2F",   x"F7",   x"DF",   x"A7",   x"8F", 
  x"D4",   x"FC",   x"84",   x"AC",   x"74",   x"5C",   x"24",   x"0C", 
  x"DB",   x"F3",   x"8B",   x"A3",   x"7B",   x"53",   x"2B",   x"03", 
  x"58",   x"70",   x"08",   x"20",   x"F8",   x"D0",   x"A8",   x"80", 
  x"1E",   x"36",   x"4E",   x"66",   x"BE",   x"96",   x"EE",   x"C6", 
  x"9D",   x"B5",   x"CD",   x"E5",   x"3D",   x"15",   x"6D",   x"45", 
  x"E7",   x"CF",   x"B7",   x"9F",   x"47",   x"6F",   x"17",   x"3F", 
  x"64",   x"4C",   x"34",   x"1C",   x"C4",   x"EC",   x"94",   x"BC", 
  x"22",   x"0A",   x"72",   x"5A",   x"82",   x"AA",   x"D2",   x"FA", 
  x"A1",   x"89",   x"F1",   x"D9",   x"01",   x"29",   x"51",   x"79", 
  x"AE",   x"86",   x"FE",   x"D6",   x"0E",   x"26",   x"5E",   x"76", 
  x"2D",   x"05",   x"7D",   x"55",   x"8D",   x"A5",   x"DD",   x"F5", 
  x"6B",   x"43",   x"3B",   x"13",   x"CB",   x"E3",   x"9B",   x"B3", 
  x"E8",   x"C0",   x"B8",   x"90",   x"48",   x"60",   x"18",   x"30", 
  x"75",   x"5D",   x"25",   x"0D",   x"D5",   x"FD",   x"85",   x"AD", 
  x"F6",   x"DE",   x"A6",   x"8E",   x"56",   x"7E",   x"06",   x"2E", 
  x"B0",   x"98",   x"E0",   x"C8",   x"10",   x"38",   x"40",   x"68", 
  x"33",   x"1B",   x"63",   x"4B",   x"93",   x"BB",   x"C3",   x"EB", 
  x"3C",   x"14",   x"6C",   x"44",   x"9C",   x"B4",   x"CC",   x"E4", 
  x"BF",   x"97",   x"EF",   x"C7",   x"1F",   x"37",   x"4F",   x"67", 
  x"F9",   x"D1",   x"A9",   x"81",   x"59",   x"71",   x"09",   x"21", 
  x"7A",   x"52",   x"2A",   x"02",   x"DA",   x"F2",   x"8A",   x"A2", 
  x"00",   x"29",   x"52",   x"7B",   x"A4",   x"8D",   x"F6",   x"DF", 
  x"8B",   x"A2",   x"D9",   x"F0",   x"2F",   x"06",   x"7D",   x"54", 
  x"D5",   x"FC",   x"87",   x"AE",   x"71",   x"58",   x"23",   x"0A", 
  x"5E",   x"77",   x"0C",   x"25",   x"FA",   x"D3",   x"A8",   x"81", 
  x"69",   x"40",   x"3B",   x"12",   x"CD",   x"E4",   x"9F",   x"B6", 
  x"E2",   x"CB",   x"B0",   x"99",   x"46",   x"6F",   x"14",   x"3D", 
  x"BC",   x"95",   x"EE",   x"C7",   x"18",   x"31",   x"4A",   x"63", 
  x"37",   x"1E",   x"65",   x"4C",   x"93",   x"BA",   x"C1",   x"E8", 
  x"D2",   x"FB",   x"80",   x"A9",   x"76",   x"5F",   x"24",   x"0D", 
  x"59",   x"70",   x"0B",   x"22",   x"FD",   x"D4",   x"AF",   x"86", 
  x"07",   x"2E",   x"55",   x"7C",   x"A3",   x"8A",   x"F1",   x"D8", 
  x"8C",   x"A5",   x"DE",   x"F7",   x"28",   x"01",   x"7A",   x"53", 
  x"BB",   x"92",   x"E9",   x"C0",   x"1F",   x"36",   x"4D",   x"64", 
  x"30",   x"19",   x"62",   x"4B",   x"94",   x"BD",   x"C6",   x"EF", 
  x"6E",   x"47",   x"3C",   x"15",   x"CA",   x"E3",   x"98",   x"B1", 
  x"E5",   x"CC",   x"B7",   x"9E",   x"41",   x"68",   x"13",   x"3A", 
  x"67",   x"4E",   x"35",   x"1C",   x"C3",   x"EA",   x"91",   x"B8", 
  x"EC",   x"C5",   x"BE",   x"97",   x"48",   x"61",   x"1A",   x"33", 
  x"B2",   x"9B",   x"E0",   x"C9",   x"16",   x"3F",   x"44",   x"6D", 
  x"39",   x"10",   x"6B",   x"42",   x"9D",   x"B4",   x"CF",   x"E6", 
  x"0E",   x"27",   x"5C",   x"75",   x"AA",   x"83",   x"F8",   x"D1", 
  x"85",   x"AC",   x"D7",   x"FE",   x"21",   x"08",   x"73",   x"5A", 
  x"DB",   x"F2",   x"89",   x"A0",   x"7F",   x"56",   x"2D",   x"04", 
  x"50",   x"79",   x"02",   x"2B",   x"F4",   x"DD",   x"A6",   x"8F", 
  x"B5",   x"9C",   x"E7",   x"CE",   x"11",   x"38",   x"43",   x"6A", 
  x"3E",   x"17",   x"6C",   x"45",   x"9A",   x"B3",   x"C8",   x"E1", 
  x"60",   x"49",   x"32",   x"1B",   x"C4",   x"ED",   x"96",   x"BF", 
  x"EB",   x"C2",   x"B9",   x"90",   x"4F",   x"66",   x"1D",   x"34", 
  x"DC",   x"F5",   x"8E",   x"A7",   x"78",   x"51",   x"2A",   x"03", 
  x"57",   x"7E",   x"05",   x"2C",   x"F3",   x"DA",   x"A1",   x"88", 
  x"09",   x"20",   x"5B",   x"72",   x"AD",   x"84",   x"FF",   x"D6", 
  x"82",   x"AB",   x"D0",   x"F9",   x"26",   x"0F",   x"74",   x"5D", 
  x"00",   x"2A",   x"54",   x"7E",   x"A8",   x"82",   x"FC",   x"D6", 
  x"93",   x"B9",   x"C7",   x"ED",   x"3B",   x"11",   x"6F",   x"45", 
  x"E5",   x"CF",   x"B1",   x"9B",   x"4D",   x"67",   x"19",   x"33", 
  x"76",   x"5C",   x"22",   x"08",   x"DE",   x"F4",   x"8A",   x"A0", 
  x"09",   x"23",   x"5D",   x"77",   x"A1",   x"8B",   x"F5",   x"DF", 
  x"9A",   x"B0",   x"CE",   x"E4",   x"32",   x"18",   x"66",   x"4C", 
  x"EC",   x"C6",   x"B8",   x"92",   x"44",   x"6E",   x"10",   x"3A", 
  x"7F",   x"55",   x"2B",   x"01",   x"D7",   x"FD",   x"83",   x"A9", 
  x"12",   x"38",   x"46",   x"6C",   x"BA",   x"90",   x"EE",   x"C4", 
  x"81",   x"AB",   x"D5",   x"FF",   x"29",   x"03",   x"7D",   x"57", 
  x"F7",   x"DD",   x"A3",   x"89",   x"5F",   x"75",   x"0B",   x"21", 
  x"64",   x"4E",   x"30",   x"1A",   x"CC",   x"E6",   x"98",   x"B2", 
  x"1B",   x"31",   x"4F",   x"65",   x"B3",   x"99",   x"E7",   x"CD", 
  x"88",   x"A2",   x"DC",   x"F6",   x"20",   x"0A",   x"74",   x"5E", 
  x"FE",   x"D4",   x"AA",   x"80",   x"56",   x"7C",   x"02",   x"28", 
  x"6D",   x"47",   x"39",   x"13",   x"C5",   x"EF",   x"91",   x"BB", 
  x"24",   x"0E",   x"70",   x"5A",   x"8C",   x"A6",   x"D8",   x"F2", 
  x"B7",   x"9D",   x"E3",   x"C9",   x"1F",   x"35",   x"4B",   x"61", 
  x"C1",   x"EB",   x"95",   x"BF",   x"69",   x"43",   x"3D",   x"17", 
  x"52",   x"78",   x"06",   x"2C",   x"FA",   x"D0",   x"AE",   x"84", 
  x"2D",   x"07",   x"79",   x"53",   x"85",   x"AF",   x"D1",   x"FB", 
  x"BE",   x"94",   x"EA",   x"C0",   x"16",   x"3C",   x"42",   x"68", 
  x"C8",   x"E2",   x"9C",   x"B6",   x"60",   x"4A",   x"34",   x"1E", 
  x"5B",   x"71",   x"0F",   x"25",   x"F3",   x"D9",   x"A7",   x"8D", 
  x"36",   x"1C",   x"62",   x"48",   x"9E",   x"B4",   x"CA",   x"E0", 
  x"A5",   x"8F",   x"F1",   x"DB",   x"0D",   x"27",   x"59",   x"73", 
  x"D3",   x"F9",   x"87",   x"AD",   x"7B",   x"51",   x"2F",   x"05", 
  x"40",   x"6A",   x"14",   x"3E",   x"E8",   x"C2",   x"BC",   x"96", 
  x"3F",   x"15",   x"6B",   x"41",   x"97",   x"BD",   x"C3",   x"E9", 
  x"AC",   x"86",   x"F8",   x"D2",   x"04",   x"2E",   x"50",   x"7A", 
  x"DA",   x"F0",   x"8E",   x"A4",   x"72",   x"58",   x"26",   x"0C", 
  x"49",   x"63",   x"1D",   x"37",   x"E1",   x"CB",   x"B5",   x"9F", 
  x"00",   x"2B",   x"56",   x"7D",   x"AC",   x"87",   x"FA",   x"D1", 
  x"9B",   x"B0",   x"CD",   x"E6",   x"37",   x"1C",   x"61",   x"4A", 
  x"F5",   x"DE",   x"A3",   x"88",   x"59",   x"72",   x"0F",   x"24", 
  x"6E",   x"45",   x"38",   x"13",   x"C2",   x"E9",   x"94",   x"BF", 
  x"29",   x"02",   x"7F",   x"54",   x"85",   x"AE",   x"D3",   x"F8", 
  x"B2",   x"99",   x"E4",   x"CF",   x"1E",   x"35",   x"48",   x"63", 
  x"DC",   x"F7",   x"8A",   x"A1",   x"70",   x"5B",   x"26",   x"0D", 
  x"47",   x"6C",   x"11",   x"3A",   x"EB",   x"C0",   x"BD",   x"96", 
  x"52",   x"79",   x"04",   x"2F",   x"FE",   x"D5",   x"A8",   x"83", 
  x"C9",   x"E2",   x"9F",   x"B4",   x"65",   x"4E",   x"33",   x"18", 
  x"A7",   x"8C",   x"F1",   x"DA",   x"0B",   x"20",   x"5D",   x"76", 
  x"3C",   x"17",   x"6A",   x"41",   x"90",   x"BB",   x"C6",   x"ED", 
  x"7B",   x"50",   x"2D",   x"06",   x"D7",   x"FC",   x"81",   x"AA", 
  x"E0",   x"CB",   x"B6",   x"9D",   x"4C",   x"67",   x"1A",   x"31", 
  x"8E",   x"A5",   x"D8",   x"F3",   x"22",   x"09",   x"74",   x"5F", 
  x"15",   x"3E",   x"43",   x"68",   x"B9",   x"92",   x"EF",   x"C4", 
  x"A4",   x"8F",   x"F2",   x"D9",   x"08",   x"23",   x"5E",   x"75", 
  x"3F",   x"14",   x"69",   x"42",   x"93",   x"B8",   x"C5",   x"EE", 
  x"51",   x"7A",   x"07",   x"2C",   x"FD",   x"D6",   x"AB",   x"80", 
  x"CA",   x"E1",   x"9C",   x"B7",   x"66",   x"4D",   x"30",   x"1B", 
  x"8D",   x"A6",   x"DB",   x"F0",   x"21",   x"0A",   x"77",   x"5C", 
  x"16",   x"3D",   x"40",   x"6B",   x"BA",   x"91",   x"EC",   x"C7", 
  x"78",   x"53",   x"2E",   x"05",   x"D4",   x"FF",   x"82",   x"A9", 
  x"E3",   x"C8",   x"B5",   x"9E",   x"4F",   x"64",   x"19",   x"32", 
  x"F6",   x"DD",   x"A0",   x"8B",   x"5A",   x"71",   x"0C",   x"27", 
  x"6D",   x"46",   x"3B",   x"10",   x"C1",   x"EA",   x"97",   x"BC", 
  x"03",   x"28",   x"55",   x"7E",   x"AF",   x"84",   x"F9",   x"D2", 
  x"98",   x"B3",   x"CE",   x"E5",   x"34",   x"1F",   x"62",   x"49", 
  x"DF",   x"F4",   x"89",   x"A2",   x"73",   x"58",   x"25",   x"0E", 
  x"44",   x"6F",   x"12",   x"39",   x"E8",   x"C3",   x"BE",   x"95", 
  x"2A",   x"01",   x"7C",   x"57",   x"86",   x"AD",   x"D0",   x"FB", 
  x"B1",   x"9A",   x"E7",   x"CC",   x"1D",   x"36",   x"4B",   x"60", 
  x"00",   x"2C",   x"58",   x"74",   x"B0",   x"9C",   x"E8",   x"C4", 
  x"A3",   x"8F",   x"FB",   x"D7",   x"13",   x"3F",   x"4B",   x"67", 
  x"85",   x"A9",   x"DD",   x"F1",   x"35",   x"19",   x"6D",   x"41", 
  x"26",   x"0A",   x"7E",   x"52",   x"96",   x"BA",   x"CE",   x"E2", 
  x"C9",   x"E5",   x"91",   x"BD",   x"79",   x"55",   x"21",   x"0D", 
  x"6A",   x"46",   x"32",   x"1E",   x"DA",   x"F6",   x"82",   x"AE", 
  x"4C",   x"60",   x"14",   x"38",   x"FC",   x"D0",   x"A4",   x"88", 
  x"EF",   x"C3",   x"B7",   x"9B",   x"5F",   x"73",   x"07",   x"2B", 
  x"51",   x"7D",   x"09",   x"25",   x"E1",   x"CD",   x"B9",   x"95", 
  x"F2",   x"DE",   x"AA",   x"86",   x"42",   x"6E",   x"1A",   x"36", 
  x"D4",   x"F8",   x"8C",   x"A0",   x"64",   x"48",   x"3C",   x"10", 
  x"77",   x"5B",   x"2F",   x"03",   x"C7",   x"EB",   x"9F",   x"B3", 
  x"98",   x"B4",   x"C0",   x"EC",   x"28",   x"04",   x"70",   x"5C", 
  x"3B",   x"17",   x"63",   x"4F",   x"8B",   x"A7",   x"D3",   x"FF", 
  x"1D",   x"31",   x"45",   x"69",   x"AD",   x"81",   x"F5",   x"D9", 
  x"BE",   x"92",   x"E6",   x"CA",   x"0E",   x"22",   x"56",   x"7A", 
  x"A2",   x"8E",   x"FA",   x"D6",   x"12",   x"3E",   x"4A",   x"66", 
  x"01",   x"2D",   x"59",   x"75",   x"B1",   x"9D",   x"E9",   x"C5", 
  x"27",   x"0B",   x"7F",   x"53",   x"97",   x"BB",   x"CF",   x"E3", 
  x"84",   x"A8",   x"DC",   x"F0",   x"34",   x"18",   x"6C",   x"40", 
  x"6B",   x"47",   x"33",   x"1F",   x"DB",   x"F7",   x"83",   x"AF", 
  x"C8",   x"E4",   x"90",   x"BC",   x"78",   x"54",   x"20",   x"0C", 
  x"EE",   x"C2",   x"B6",   x"9A",   x"5E",   x"72",   x"06",   x"2A", 
  x"4D",   x"61",   x"15",   x"39",   x"FD",   x"D1",   x"A5",   x"89", 
  x"F3",   x"DF",   x"AB",   x"87",   x"43",   x"6F",   x"1B",   x"37", 
  x"50",   x"7C",   x"08",   x"24",   x"E0",   x"CC",   x"B8",   x"94", 
  x"76",   x"5A",   x"2E",   x"02",   x"C6",   x"EA",   x"9E",   x"B2", 
  x"D5",   x"F9",   x"8D",   x"A1",   x"65",   x"49",   x"3D",   x"11", 
  x"3A",   x"16",   x"62",   x"4E",   x"8A",   x"A6",   x"D2",   x"FE", 
  x"99",   x"B5",   x"C1",   x"ED",   x"29",   x"05",   x"71",   x"5D", 
  x"BF",   x"93",   x"E7",   x"CB",   x"0F",   x"23",   x"57",   x"7B", 
  x"1C",   x"30",   x"44",   x"68",   x"AC",   x"80",   x"F4",   x"D8", 
  x"00",   x"2D",   x"5A",   x"77",   x"B4",   x"99",   x"EE",   x"C3", 
  x"AB",   x"86",   x"F1",   x"DC",   x"1F",   x"32",   x"45",   x"68", 
  x"95",   x"B8",   x"CF",   x"E2",   x"21",   x"0C",   x"7B",   x"56", 
  x"3E",   x"13",   x"64",   x"49",   x"8A",   x"A7",   x"D0",   x"FD", 
  x"E9",   x"C4",   x"B3",   x"9E",   x"5D",   x"70",   x"07",   x"2A", 
  x"42",   x"6F",   x"18",   x"35",   x"F6",   x"DB",   x"AC",   x"81", 
  x"7C",   x"51",   x"26",   x"0B",   x"C8",   x"E5",   x"92",   x"BF", 
  x"D7",   x"FA",   x"8D",   x"A0",   x"63",   x"4E",   x"39",   x"14", 
  x"11",   x"3C",   x"4B",   x"66",   x"A5",   x"88",   x"FF",   x"D2", 
  x"BA",   x"97",   x"E0",   x"CD",   x"0E",   x"23",   x"54",   x"79", 
  x"84",   x"A9",   x"DE",   x"F3",   x"30",   x"1D",   x"6A",   x"47", 
  x"2F",   x"02",   x"75",   x"58",   x"9B",   x"B6",   x"C1",   x"EC", 
  x"F8",   x"D5",   x"A2",   x"8F",   x"4C",   x"61",   x"16",   x"3B", 
  x"53",   x"7E",   x"09",   x"24",   x"E7",   x"CA",   x"BD",   x"90", 
  x"6D",   x"40",   x"37",   x"1A",   x"D9",   x"F4",   x"83",   x"AE", 
  x"C6",   x"EB",   x"9C",   x"B1",   x"72",   x"5F",   x"28",   x"05", 
  x"22",   x"0F",   x"78",   x"55",   x"96",   x"BB",   x"CC",   x"E1", 
  x"89",   x"A4",   x"D3",   x"FE",   x"3D",   x"10",   x"67",   x"4A", 
  x"B7",   x"9A",   x"ED",   x"C0",   x"03",   x"2E",   x"59",   x"74", 
  x"1C",   x"31",   x"46",   x"6B",   x"A8",   x"85",   x"F2",   x"DF", 
  x"CB",   x"E6",   x"91",   x"BC",   x"7F",   x"52",   x"25",   x"08", 
  x"60",   x"4D",   x"3A",   x"17",   x"D4",   x"F9",   x"8E",   x"A3", 
  x"5E",   x"73",   x"04",   x"29",   x"EA",   x"C7",   x"B0",   x"9D", 
  x"F5",   x"D8",   x"AF",   x"82",   x"41",   x"6C",   x"1B",   x"36", 
  x"33",   x"1E",   x"69",   x"44",   x"87",   x"AA",   x"DD",   x"F0", 
  x"98",   x"B5",   x"C2",   x"EF",   x"2C",   x"01",   x"76",   x"5B", 
  x"A6",   x"8B",   x"FC",   x"D1",   x"12",   x"3F",   x"48",   x"65", 
  x"0D",   x"20",   x"57",   x"7A",   x"B9",   x"94",   x"E3",   x"CE", 
  x"DA",   x"F7",   x"80",   x"AD",   x"6E",   x"43",   x"34",   x"19", 
  x"71",   x"5C",   x"2B",   x"06",   x"C5",   x"E8",   x"9F",   x"B2", 
  x"4F",   x"62",   x"15",   x"38",   x"FB",   x"D6",   x"A1",   x"8C", 
  x"E4",   x"C9",   x"BE",   x"93",   x"50",   x"7D",   x"0A",   x"27", 
  x"00",   x"2E",   x"5C",   x"72",   x"B8",   x"96",   x"E4",   x"CA", 
  x"B3",   x"9D",   x"EF",   x"C1",   x"0B",   x"25",   x"57",   x"79", 
  x"A5",   x"8B",   x"F9",   x"D7",   x"1D",   x"33",   x"41",   x"6F", 
  x"16",   x"38",   x"4A",   x"64",   x"AE",   x"80",   x"F2",   x"DC", 
  x"89",   x"A7",   x"D5",   x"FB",   x"31",   x"1F",   x"6D",   x"43", 
  x"3A",   x"14",   x"66",   x"48",   x"82",   x"AC",   x"DE",   x"F0", 
  x"2C",   x"02",   x"70",   x"5E",   x"94",   x"BA",   x"C8",   x"E6", 
  x"9F",   x"B1",   x"C3",   x"ED",   x"27",   x"09",   x"7B",   x"55", 
  x"D1",   x"FF",   x"8D",   x"A3",   x"69",   x"47",   x"35",   x"1B", 
  x"62",   x"4C",   x"3E",   x"10",   x"DA",   x"F4",   x"86",   x"A8", 
  x"74",   x"5A",   x"28",   x"06",   x"CC",   x"E2",   x"90",   x"BE", 
  x"C7",   x"E9",   x"9B",   x"B5",   x"7F",   x"51",   x"23",   x"0D", 
  x"58",   x"76",   x"04",   x"2A",   x"E0",   x"CE",   x"BC",   x"92", 
  x"EB",   x"C5",   x"B7",   x"99",   x"53",   x"7D",   x"0F",   x"21", 
  x"FD",   x"D3",   x"A1",   x"8F",   x"45",   x"6B",   x"19",   x"37", 
  x"4E",   x"60",   x"12",   x"3C",   x"F6",   x"D8",   x"AA",   x"84", 
  x"61",   x"4F",   x"3D",   x"13",   x"D9",   x"F7",   x"85",   x"AB", 
  x"D2",   x"FC",   x"8E",   x"A0",   x"6A",   x"44",   x"36",   x"18", 
  x"C4",   x"EA",   x"98",   x"B6",   x"7C",   x"52",   x"20",   x"0E", 
  x"77",   x"59",   x"2B",   x"05",   x"CF",   x"E1",   x"93",   x"BD", 
  x"E8",   x"C6",   x"B4",   x"9A",   x"50",   x"7E",   x"0C",   x"22", 
  x"5B",   x"75",   x"07",   x"29",   x"E3",   x"CD",   x"BF",   x"91", 
  x"4D",   x"63",   x"11",   x"3F",   x"F5",   x"DB",   x"A9",   x"87", 
  x"FE",   x"D0",   x"A2",   x"8C",   x"46",   x"68",   x"1A",   x"34", 
  x"B0",   x"9E",   x"EC",   x"C2",   x"08",   x"26",   x"54",   x"7A", 
  x"03",   x"2D",   x"5F",   x"71",   x"BB",   x"95",   x"E7",   x"C9", 
  x"15",   x"3B",   x"49",   x"67",   x"AD",   x"83",   x"F1",   x"DF", 
  x"A6",   x"88",   x"FA",   x"D4",   x"1E",   x"30",   x"42",   x"6C", 
  x"39",   x"17",   x"65",   x"4B",   x"81",   x"AF",   x"DD",   x"F3", 
  x"8A",   x"A4",   x"D6",   x"F8",   x"32",   x"1C",   x"6E",   x"40", 
  x"9C",   x"B2",   x"C0",   x"EE",   x"24",   x"0A",   x"78",   x"56", 
  x"2F",   x"01",   x"73",   x"5D",   x"97",   x"B9",   x"CB",   x"E5", 
  x"00",   x"2F",   x"5E",   x"71",   x"BC",   x"93",   x"E2",   x"CD", 
  x"BB",   x"94",   x"E5",   x"CA",   x"07",   x"28",   x"59",   x"76", 
  x"B5",   x"9A",   x"EB",   x"C4",   x"09",   x"26",   x"57",   x"78", 
  x"0E",   x"21",   x"50",   x"7F",   x"B2",   x"9D",   x"EC",   x"C3", 
  x"A9",   x"86",   x"F7",   x"D8",   x"15",   x"3A",   x"4B",   x"64", 
  x"12",   x"3D",   x"4C",   x"63",   x"AE",   x"81",   x"F0",   x"DF", 
  x"1C",   x"33",   x"42",   x"6D",   x"A0",   x"8F",   x"FE",   x"D1", 
  x"A7",   x"88",   x"F9",   x"D6",   x"1B",   x"34",   x"45",   x"6A", 
  x"91",   x"BE",   x"CF",   x"E0",   x"2D",   x"02",   x"73",   x"5C", 
  x"2A",   x"05",   x"74",   x"5B",   x"96",   x"B9",   x"C8",   x"E7", 
  x"24",   x"0B",   x"7A",   x"55",   x"98",   x"B7",   x"C6",   x"E9", 
  x"9F",   x"B0",   x"C1",   x"EE",   x"23",   x"0C",   x"7D",   x"52", 
  x"38",   x"17",   x"66",   x"49",   x"84",   x"AB",   x"DA",   x"F5", 
  x"83",   x"AC",   x"DD",   x"F2",   x"3F",   x"10",   x"61",   x"4E", 
  x"8D",   x"A2",   x"D3",   x"FC",   x"31",   x"1E",   x"6F",   x"40", 
  x"36",   x"19",   x"68",   x"47",   x"8A",   x"A5",   x"D4",   x"FB", 
  x"E1",   x"CE",   x"BF",   x"90",   x"5D",   x"72",   x"03",   x"2C", 
  x"5A",   x"75",   x"04",   x"2B",   x"E6",   x"C9",   x"B8",   x"97", 
  x"54",   x"7B",   x"0A",   x"25",   x"E8",   x"C7",   x"B6",   x"99", 
  x"EF",   x"C0",   x"B1",   x"9E",   x"53",   x"7C",   x"0D",   x"22", 
  x"48",   x"67",   x"16",   x"39",   x"F4",   x"DB",   x"AA",   x"85", 
  x"F3",   x"DC",   x"AD",   x"82",   x"4F",   x"60",   x"11",   x"3E", 
  x"FD",   x"D2",   x"A3",   x"8C",   x"41",   x"6E",   x"1F",   x"30", 
  x"46",   x"69",   x"18",   x"37",   x"FA",   x"D5",   x"A4",   x"8B", 
  x"70",   x"5F",   x"2E",   x"01",   x"CC",   x"E3",   x"92",   x"BD", 
  x"CB",   x"E4",   x"95",   x"BA",   x"77",   x"58",   x"29",   x"06", 
  x"C5",   x"EA",   x"9B",   x"B4",   x"79",   x"56",   x"27",   x"08", 
  x"7E",   x"51",   x"20",   x"0F",   x"C2",   x"ED",   x"9C",   x"B3", 
  x"D9",   x"F6",   x"87",   x"A8",   x"65",   x"4A",   x"3B",   x"14", 
  x"62",   x"4D",   x"3C",   x"13",   x"DE",   x"F1",   x"80",   x"AF", 
  x"6C",   x"43",   x"32",   x"1D",   x"D0",   x"FF",   x"8E",   x"A1", 
  x"D7",   x"F8",   x"89",   x"A6",   x"6B",   x"44",   x"35",   x"1A", 
  x"00",   x"30",   x"60",   x"50",   x"C0",   x"F0",   x"A0",   x"90", 
  x"43",   x"73",   x"23",   x"13",   x"83",   x"B3",   x"E3",   x"D3", 
  x"86",   x"B6",   x"E6",   x"D6",   x"46",   x"76",   x"26",   x"16", 
  x"C5",   x"F5",   x"A5",   x"95",   x"05",   x"35",   x"65",   x"55", 
  x"CF",   x"FF",   x"AF",   x"9F",   x"0F",   x"3F",   x"6F",   x"5F", 
  x"8C",   x"BC",   x"EC",   x"DC",   x"4C",   x"7C",   x"2C",   x"1C", 
  x"49",   x"79",   x"29",   x"19",   x"89",   x"B9",   x"E9",   x"D9", 
  x"0A",   x"3A",   x"6A",   x"5A",   x"CA",   x"FA",   x"AA",   x"9A", 
  x"5D",   x"6D",   x"3D",   x"0D",   x"9D",   x"AD",   x"FD",   x"CD", 
  x"1E",   x"2E",   x"7E",   x"4E",   x"DE",   x"EE",   x"BE",   x"8E", 
  x"DB",   x"EB",   x"BB",   x"8B",   x"1B",   x"2B",   x"7B",   x"4B", 
  x"98",   x"A8",   x"F8",   x"C8",   x"58",   x"68",   x"38",   x"08", 
  x"92",   x"A2",   x"F2",   x"C2",   x"52",   x"62",   x"32",   x"02", 
  x"D1",   x"E1",   x"B1",   x"81",   x"11",   x"21",   x"71",   x"41", 
  x"14",   x"24",   x"74",   x"44",   x"D4",   x"E4",   x"B4",   x"84", 
  x"57",   x"67",   x"37",   x"07",   x"97",   x"A7",   x"F7",   x"C7", 
  x"BA",   x"8A",   x"DA",   x"EA",   x"7A",   x"4A",   x"1A",   x"2A", 
  x"F9",   x"C9",   x"99",   x"A9",   x"39",   x"09",   x"59",   x"69", 
  x"3C",   x"0C",   x"5C",   x"6C",   x"FC",   x"CC",   x"9C",   x"AC", 
  x"7F",   x"4F",   x"1F",   x"2F",   x"BF",   x"8F",   x"DF",   x"EF", 
  x"75",   x"45",   x"15",   x"25",   x"B5",   x"85",   x"D5",   x"E5", 
  x"36",   x"06",   x"56",   x"66",   x"F6",   x"C6",   x"96",   x"A6", 
  x"F3",   x"C3",   x"93",   x"A3",   x"33",   x"03",   x"53",   x"63", 
  x"B0",   x"80",   x"D0",   x"E0",   x"70",   x"40",   x"10",   x"20", 
  x"E7",   x"D7",   x"87",   x"B7",   x"27",   x"17",   x"47",   x"77", 
  x"A4",   x"94",   x"C4",   x"F4",   x"64",   x"54",   x"04",   x"34", 
  x"61",   x"51",   x"01",   x"31",   x"A1",   x"91",   x"C1",   x"F1", 
  x"22",   x"12",   x"42",   x"72",   x"E2",   x"D2",   x"82",   x"B2", 
  x"28",   x"18",   x"48",   x"78",   x"E8",   x"D8",   x"88",   x"B8", 
  x"6B",   x"5B",   x"0B",   x"3B",   x"AB",   x"9B",   x"CB",   x"FB", 
  x"AE",   x"9E",   x"CE",   x"FE",   x"6E",   x"5E",   x"0E",   x"3E", 
  x"ED",   x"DD",   x"8D",   x"BD",   x"2D",   x"1D",   x"4D",   x"7D", 
  x"00",   x"31",   x"62",   x"53",   x"C4",   x"F5",   x"A6",   x"97", 
  x"4B",   x"7A",   x"29",   x"18",   x"8F",   x"BE",   x"ED",   x"DC", 
  x"96",   x"A7",   x"F4",   x"C5",   x"52",   x"63",   x"30",   x"01", 
  x"DD",   x"EC",   x"BF",   x"8E",   x"19",   x"28",   x"7B",   x"4A", 
  x"EF",   x"DE",   x"8D",   x"BC",   x"2B",   x"1A",   x"49",   x"78", 
  x"A4",   x"95",   x"C6",   x"F7",   x"60",   x"51",   x"02",   x"33", 
  x"79",   x"48",   x"1B",   x"2A",   x"BD",   x"8C",   x"DF",   x"EE", 
  x"32",   x"03",   x"50",   x"61",   x"F6",   x"C7",   x"94",   x"A5", 
  x"1D",   x"2C",   x"7F",   x"4E",   x"D9",   x"E8",   x"BB",   x"8A", 
  x"56",   x"67",   x"34",   x"05",   x"92",   x"A3",   x"F0",   x"C1", 
  x"8B",   x"BA",   x"E9",   x"D8",   x"4F",   x"7E",   x"2D",   x"1C", 
  x"C0",   x"F1",   x"A2",   x"93",   x"04",   x"35",   x"66",   x"57", 
  x"F2",   x"C3",   x"90",   x"A1",   x"36",   x"07",   x"54",   x"65", 
  x"B9",   x"88",   x"DB",   x"EA",   x"7D",   x"4C",   x"1F",   x"2E", 
  x"64",   x"55",   x"06",   x"37",   x"A0",   x"91",   x"C2",   x"F3", 
  x"2F",   x"1E",   x"4D",   x"7C",   x"EB",   x"DA",   x"89",   x"B8", 
  x"3A",   x"0B",   x"58",   x"69",   x"FE",   x"CF",   x"9C",   x"AD", 
  x"71",   x"40",   x"13",   x"22",   x"B5",   x"84",   x"D7",   x"E6", 
  x"AC",   x"9D",   x"CE",   x"FF",   x"68",   x"59",   x"0A",   x"3B", 
  x"E7",   x"D6",   x"85",   x"B4",   x"23",   x"12",   x"41",   x"70", 
  x"D5",   x"E4",   x"B7",   x"86",   x"11",   x"20",   x"73",   x"42", 
  x"9E",   x"AF",   x"FC",   x"CD",   x"5A",   x"6B",   x"38",   x"09", 
  x"43",   x"72",   x"21",   x"10",   x"87",   x"B6",   x"E5",   x"D4", 
  x"08",   x"39",   x"6A",   x"5B",   x"CC",   x"FD",   x"AE",   x"9F", 
  x"27",   x"16",   x"45",   x"74",   x"E3",   x"D2",   x"81",   x"B0", 
  x"6C",   x"5D",   x"0E",   x"3F",   x"A8",   x"99",   x"CA",   x"FB", 
  x"B1",   x"80",   x"D3",   x"E2",   x"75",   x"44",   x"17",   x"26", 
  x"FA",   x"CB",   x"98",   x"A9",   x"3E",   x"0F",   x"5C",   x"6D", 
  x"C8",   x"F9",   x"AA",   x"9B",   x"0C",   x"3D",   x"6E",   x"5F", 
  x"83",   x"B2",   x"E1",   x"D0",   x"47",   x"76",   x"25",   x"14", 
  x"5E",   x"6F",   x"3C",   x"0D",   x"9A",   x"AB",   x"F8",   x"C9", 
  x"15",   x"24",   x"77",   x"46",   x"D1",   x"E0",   x"B3",   x"82", 
  x"00",   x"32",   x"64",   x"56",   x"C8",   x"FA",   x"AC",   x"9E", 
  x"53",   x"61",   x"37",   x"05",   x"9B",   x"A9",   x"FF",   x"CD", 
  x"A6",   x"94",   x"C2",   x"F0",   x"6E",   x"5C",   x"0A",   x"38", 
  x"F5",   x"C7",   x"91",   x"A3",   x"3D",   x"0F",   x"59",   x"6B", 
  x"8F",   x"BD",   x"EB",   x"D9",   x"47",   x"75",   x"23",   x"11", 
  x"DC",   x"EE",   x"B8",   x"8A",   x"14",   x"26",   x"70",   x"42", 
  x"29",   x"1B",   x"4D",   x"7F",   x"E1",   x"D3",   x"85",   x"B7", 
  x"7A",   x"48",   x"1E",   x"2C",   x"B2",   x"80",   x"D6",   x"E4", 
  x"DD",   x"EF",   x"B9",   x"8B",   x"15",   x"27",   x"71",   x"43", 
  x"8E",   x"BC",   x"EA",   x"D8",   x"46",   x"74",   x"22",   x"10", 
  x"7B",   x"49",   x"1F",   x"2D",   x"B3",   x"81",   x"D7",   x"E5", 
  x"28",   x"1A",   x"4C",   x"7E",   x"E0",   x"D2",   x"84",   x"B6", 
  x"52",   x"60",   x"36",   x"04",   x"9A",   x"A8",   x"FE",   x"CC", 
  x"01",   x"33",   x"65",   x"57",   x"C9",   x"FB",   x"AD",   x"9F", 
  x"F4",   x"C6",   x"90",   x"A2",   x"3C",   x"0E",   x"58",   x"6A", 
  x"A7",   x"95",   x"C3",   x"F1",   x"6F",   x"5D",   x"0B",   x"39", 
  x"79",   x"4B",   x"1D",   x"2F",   x"B1",   x"83",   x"D5",   x"E7", 
  x"2A",   x"18",   x"4E",   x"7C",   x"E2",   x"D0",   x"86",   x"B4", 
  x"DF",   x"ED",   x"BB",   x"89",   x"17",   x"25",   x"73",   x"41", 
  x"8C",   x"BE",   x"E8",   x"DA",   x"44",   x"76",   x"20",   x"12", 
  x"F6",   x"C4",   x"92",   x"A0",   x"3E",   x"0C",   x"5A",   x"68", 
  x"A5",   x"97",   x"C1",   x"F3",   x"6D",   x"5F",   x"09",   x"3B", 
  x"50",   x"62",   x"34",   x"06",   x"98",   x"AA",   x"FC",   x"CE", 
  x"03",   x"31",   x"67",   x"55",   x"CB",   x"F9",   x"AF",   x"9D", 
  x"A4",   x"96",   x"C0",   x"F2",   x"6C",   x"5E",   x"08",   x"3A", 
  x"F7",   x"C5",   x"93",   x"A1",   x"3F",   x"0D",   x"5B",   x"69", 
  x"02",   x"30",   x"66",   x"54",   x"CA",   x"F8",   x"AE",   x"9C", 
  x"51",   x"63",   x"35",   x"07",   x"99",   x"AB",   x"FD",   x"CF", 
  x"2B",   x"19",   x"4F",   x"7D",   x"E3",   x"D1",   x"87",   x"B5", 
  x"78",   x"4A",   x"1C",   x"2E",   x"B0",   x"82",   x"D4",   x"E6", 
  x"8D",   x"BF",   x"E9",   x"DB",   x"45",   x"77",   x"21",   x"13", 
  x"DE",   x"EC",   x"BA",   x"88",   x"16",   x"24",   x"72",   x"40", 
  x"00",   x"33",   x"66",   x"55",   x"CC",   x"FF",   x"AA",   x"99", 
  x"5B",   x"68",   x"3D",   x"0E",   x"97",   x"A4",   x"F1",   x"C2", 
  x"B6",   x"85",   x"D0",   x"E3",   x"7A",   x"49",   x"1C",   x"2F", 
  x"ED",   x"DE",   x"8B",   x"B8",   x"21",   x"12",   x"47",   x"74", 
  x"AF",   x"9C",   x"C9",   x"FA",   x"63",   x"50",   x"05",   x"36", 
  x"F4",   x"C7",   x"92",   x"A1",   x"38",   x"0B",   x"5E",   x"6D", 
  x"19",   x"2A",   x"7F",   x"4C",   x"D5",   x"E6",   x"B3",   x"80", 
  x"42",   x"71",   x"24",   x"17",   x"8E",   x"BD",   x"E8",   x"DB", 
  x"9D",   x"AE",   x"FB",   x"C8",   x"51",   x"62",   x"37",   x"04", 
  x"C6",   x"F5",   x"A0",   x"93",   x"0A",   x"39",   x"6C",   x"5F", 
  x"2B",   x"18",   x"4D",   x"7E",   x"E7",   x"D4",   x"81",   x"B2", 
  x"70",   x"43",   x"16",   x"25",   x"BC",   x"8F",   x"DA",   x"E9", 
  x"32",   x"01",   x"54",   x"67",   x"FE",   x"CD",   x"98",   x"AB", 
  x"69",   x"5A",   x"0F",   x"3C",   x"A5",   x"96",   x"C3",   x"F0", 
  x"84",   x"B7",   x"E2",   x"D1",   x"48",   x"7B",   x"2E",   x"1D", 
  x"DF",   x"EC",   x"B9",   x"8A",   x"13",   x"20",   x"75",   x"46", 
  x"F9",   x"CA",   x"9F",   x"AC",   x"35",   x"06",   x"53",   x"60", 
  x"A2",   x"91",   x"C4",   x"F7",   x"6E",   x"5D",   x"08",   x"3B", 
  x"4F",   x"7C",   x"29",   x"1A",   x"83",   x"B0",   x"E5",   x"D6", 
  x"14",   x"27",   x"72",   x"41",   x"D8",   x"EB",   x"BE",   x"8D", 
  x"56",   x"65",   x"30",   x"03",   x"9A",   x"A9",   x"FC",   x"CF", 
  x"0D",   x"3E",   x"6B",   x"58",   x"C1",   x"F2",   x"A7",   x"94", 
  x"E0",   x"D3",   x"86",   x"B5",   x"2C",   x"1F",   x"4A",   x"79", 
  x"BB",   x"88",   x"DD",   x"EE",   x"77",   x"44",   x"11",   x"22", 
  x"64",   x"57",   x"02",   x"31",   x"A8",   x"9B",   x"CE",   x"FD", 
  x"3F",   x"0C",   x"59",   x"6A",   x"F3",   x"C0",   x"95",   x"A6", 
  x"D2",   x"E1",   x"B4",   x"87",   x"1E",   x"2D",   x"78",   x"4B", 
  x"89",   x"BA",   x"EF",   x"DC",   x"45",   x"76",   x"23",   x"10", 
  x"CB",   x"F8",   x"AD",   x"9E",   x"07",   x"34",   x"61",   x"52", 
  x"90",   x"A3",   x"F6",   x"C5",   x"5C",   x"6F",   x"3A",   x"09", 
  x"7D",   x"4E",   x"1B",   x"28",   x"B1",   x"82",   x"D7",   x"E4", 
  x"26",   x"15",   x"40",   x"73",   x"EA",   x"D9",   x"8C",   x"BF", 
  x"00",   x"34",   x"68",   x"5C",   x"D0",   x"E4",   x"B8",   x"8C", 
  x"63",   x"57",   x"0B",   x"3F",   x"B3",   x"87",   x"DB",   x"EF", 
  x"C6",   x"F2",   x"AE",   x"9A",   x"16",   x"22",   x"7E",   x"4A", 
  x"A5",   x"91",   x"CD",   x"F9",   x"75",   x"41",   x"1D",   x"29", 
  x"4F",   x"7B",   x"27",   x"13",   x"9F",   x"AB",   x"F7",   x"C3", 
  x"2C",   x"18",   x"44",   x"70",   x"FC",   x"C8",   x"94",   x"A0", 
  x"89",   x"BD",   x"E1",   x"D5",   x"59",   x"6D",   x"31",   x"05", 
  x"EA",   x"DE",   x"82",   x"B6",   x"3A",   x"0E",   x"52",   x"66", 
  x"9E",   x"AA",   x"F6",   x"C2",   x"4E",   x"7A",   x"26",   x"12", 
  x"FD",   x"C9",   x"95",   x"A1",   x"2D",   x"19",   x"45",   x"71", 
  x"58",   x"6C",   x"30",   x"04",   x"88",   x"BC",   x"E0",   x"D4", 
  x"3B",   x"0F",   x"53",   x"67",   x"EB",   x"DF",   x"83",   x"B7", 
  x"D1",   x"E5",   x"B9",   x"8D",   x"01",   x"35",   x"69",   x"5D", 
  x"B2",   x"86",   x"DA",   x"EE",   x"62",   x"56",   x"0A",   x"3E", 
  x"17",   x"23",   x"7F",   x"4B",   x"C7",   x"F3",   x"AF",   x"9B", 
  x"74",   x"40",   x"1C",   x"28",   x"A4",   x"90",   x"CC",   x"F8", 
  x"FF",   x"CB",   x"97",   x"A3",   x"2F",   x"1B",   x"47",   x"73", 
  x"9C",   x"A8",   x"F4",   x"C0",   x"4C",   x"78",   x"24",   x"10", 
  x"39",   x"0D",   x"51",   x"65",   x"E9",   x"DD",   x"81",   x"B5", 
  x"5A",   x"6E",   x"32",   x"06",   x"8A",   x"BE",   x"E2",   x"D6", 
  x"B0",   x"84",   x"D8",   x"EC",   x"60",   x"54",   x"08",   x"3C", 
  x"D3",   x"E7",   x"BB",   x"8F",   x"03",   x"37",   x"6B",   x"5F", 
  x"76",   x"42",   x"1E",   x"2A",   x"A6",   x"92",   x"CE",   x"FA", 
  x"15",   x"21",   x"7D",   x"49",   x"C5",   x"F1",   x"AD",   x"99", 
  x"61",   x"55",   x"09",   x"3D",   x"B1",   x"85",   x"D9",   x"ED", 
  x"02",   x"36",   x"6A",   x"5E",   x"D2",   x"E6",   x"BA",   x"8E", 
  x"A7",   x"93",   x"CF",   x"FB",   x"77",   x"43",   x"1F",   x"2B", 
  x"C4",   x"F0",   x"AC",   x"98",   x"14",   x"20",   x"7C",   x"48", 
  x"2E",   x"1A",   x"46",   x"72",   x"FE",   x"CA",   x"96",   x"A2", 
  x"4D",   x"79",   x"25",   x"11",   x"9D",   x"A9",   x"F5",   x"C1", 
  x"E8",   x"DC",   x"80",   x"B4",   x"38",   x"0C",   x"50",   x"64", 
  x"8B",   x"BF",   x"E3",   x"D7",   x"5B",   x"6F",   x"33",   x"07", 
  x"00",   x"35",   x"6A",   x"5F",   x"D4",   x"E1",   x"BE",   x"8B", 
  x"6B",   x"5E",   x"01",   x"34",   x"BF",   x"8A",   x"D5",   x"E0", 
  x"D6",   x"E3",   x"BC",   x"89",   x"02",   x"37",   x"68",   x"5D", 
  x"BD",   x"88",   x"D7",   x"E2",   x"69",   x"5C",   x"03",   x"36", 
  x"6F",   x"5A",   x"05",   x"30",   x"BB",   x"8E",   x"D1",   x"E4", 
  x"04",   x"31",   x"6E",   x"5B",   x"D0",   x"E5",   x"BA",   x"8F", 
  x"B9",   x"8C",   x"D3",   x"E6",   x"6D",   x"58",   x"07",   x"32", 
  x"D2",   x"E7",   x"B8",   x"8D",   x"06",   x"33",   x"6C",   x"59", 
  x"DE",   x"EB",   x"B4",   x"81",   x"0A",   x"3F",   x"60",   x"55", 
  x"B5",   x"80",   x"DF",   x"EA",   x"61",   x"54",   x"0B",   x"3E", 
  x"08",   x"3D",   x"62",   x"57",   x"DC",   x"E9",   x"B6",   x"83", 
  x"63",   x"56",   x"09",   x"3C",   x"B7",   x"82",   x"DD",   x"E8", 
  x"B1",   x"84",   x"DB",   x"EE",   x"65",   x"50",   x"0F",   x"3A", 
  x"DA",   x"EF",   x"B0",   x"85",   x"0E",   x"3B",   x"64",   x"51", 
  x"67",   x"52",   x"0D",   x"38",   x"B3",   x"86",   x"D9",   x"EC", 
  x"0C",   x"39",   x"66",   x"53",   x"D8",   x"ED",   x"B2",   x"87", 
  x"7F",   x"4A",   x"15",   x"20",   x"AB",   x"9E",   x"C1",   x"F4", 
  x"14",   x"21",   x"7E",   x"4B",   x"C0",   x"F5",   x"AA",   x"9F", 
  x"A9",   x"9C",   x"C3",   x"F6",   x"7D",   x"48",   x"17",   x"22", 
  x"C2",   x"F7",   x"A8",   x"9D",   x"16",   x"23",   x"7C",   x"49", 
  x"10",   x"25",   x"7A",   x"4F",   x"C4",   x"F1",   x"AE",   x"9B", 
  x"7B",   x"4E",   x"11",   x"24",   x"AF",   x"9A",   x"C5",   x"F0", 
  x"C6",   x"F3",   x"AC",   x"99",   x"12",   x"27",   x"78",   x"4D", 
  x"AD",   x"98",   x"C7",   x"F2",   x"79",   x"4C",   x"13",   x"26", 
  x"A1",   x"94",   x"CB",   x"FE",   x"75",   x"40",   x"1F",   x"2A", 
  x"CA",   x"FF",   x"A0",   x"95",   x"1E",   x"2B",   x"74",   x"41", 
  x"77",   x"42",   x"1D",   x"28",   x"A3",   x"96",   x"C9",   x"FC", 
  x"1C",   x"29",   x"76",   x"43",   x"C8",   x"FD",   x"A2",   x"97", 
  x"CE",   x"FB",   x"A4",   x"91",   x"1A",   x"2F",   x"70",   x"45", 
  x"A5",   x"90",   x"CF",   x"FA",   x"71",   x"44",   x"1B",   x"2E", 
  x"18",   x"2D",   x"72",   x"47",   x"CC",   x"F9",   x"A6",   x"93", 
  x"73",   x"46",   x"19",   x"2C",   x"A7",   x"92",   x"CD",   x"F8", 
  x"00",   x"36",   x"6C",   x"5A",   x"D8",   x"EE",   x"B4",   x"82", 
  x"73",   x"45",   x"1F",   x"29",   x"AB",   x"9D",   x"C7",   x"F1", 
  x"E6",   x"D0",   x"8A",   x"BC",   x"3E",   x"08",   x"52",   x"64", 
  x"95",   x"A3",   x"F9",   x"CF",   x"4D",   x"7B",   x"21",   x"17", 
  x"0F",   x"39",   x"63",   x"55",   x"D7",   x"E1",   x"BB",   x"8D", 
  x"7C",   x"4A",   x"10",   x"26",   x"A4",   x"92",   x"C8",   x"FE", 
  x"E9",   x"DF",   x"85",   x"B3",   x"31",   x"07",   x"5D",   x"6B", 
  x"9A",   x"AC",   x"F6",   x"C0",   x"42",   x"74",   x"2E",   x"18", 
  x"1E",   x"28",   x"72",   x"44",   x"C6",   x"F0",   x"AA",   x"9C", 
  x"6D",   x"5B",   x"01",   x"37",   x"B5",   x"83",   x"D9",   x"EF", 
  x"F8",   x"CE",   x"94",   x"A2",   x"20",   x"16",   x"4C",   x"7A", 
  x"8B",   x"BD",   x"E7",   x"D1",   x"53",   x"65",   x"3F",   x"09", 
  x"11",   x"27",   x"7D",   x"4B",   x"C9",   x"FF",   x"A5",   x"93", 
  x"62",   x"54",   x"0E",   x"38",   x"BA",   x"8C",   x"D6",   x"E0", 
  x"F7",   x"C1",   x"9B",   x"AD",   x"2F",   x"19",   x"43",   x"75", 
  x"84",   x"B2",   x"E8",   x"DE",   x"5C",   x"6A",   x"30",   x"06", 
  x"3C",   x"0A",   x"50",   x"66",   x"E4",   x"D2",   x"88",   x"BE", 
  x"4F",   x"79",   x"23",   x"15",   x"97",   x"A1",   x"FB",   x"CD", 
  x"DA",   x"EC",   x"B6",   x"80",   x"02",   x"34",   x"6E",   x"58", 
  x"A9",   x"9F",   x"C5",   x"F3",   x"71",   x"47",   x"1D",   x"2B", 
  x"33",   x"05",   x"5F",   x"69",   x"EB",   x"DD",   x"87",   x"B1", 
  x"40",   x"76",   x"2C",   x"1A",   x"98",   x"AE",   x"F4",   x"C2", 
  x"D5",   x"E3",   x"B9",   x"8F",   x"0D",   x"3B",   x"61",   x"57", 
  x"A6",   x"90",   x"CA",   x"FC",   x"7E",   x"48",   x"12",   x"24", 
  x"22",   x"14",   x"4E",   x"78",   x"FA",   x"CC",   x"96",   x"A0", 
  x"51",   x"67",   x"3D",   x"0B",   x"89",   x"BF",   x"E5",   x"D3", 
  x"C4",   x"F2",   x"A8",   x"9E",   x"1C",   x"2A",   x"70",   x"46", 
  x"B7",   x"81",   x"DB",   x"ED",   x"6F",   x"59",   x"03",   x"35", 
  x"2D",   x"1B",   x"41",   x"77",   x"F5",   x"C3",   x"99",   x"AF", 
  x"5E",   x"68",   x"32",   x"04",   x"86",   x"B0",   x"EA",   x"DC", 
  x"CB",   x"FD",   x"A7",   x"91",   x"13",   x"25",   x"7F",   x"49", 
  x"B8",   x"8E",   x"D4",   x"E2",   x"60",   x"56",   x"0C",   x"3A", 
  x"00",   x"37",   x"6E",   x"59",   x"DC",   x"EB",   x"B2",   x"85", 
  x"7B",   x"4C",   x"15",   x"22",   x"A7",   x"90",   x"C9",   x"FE", 
  x"F6",   x"C1",   x"98",   x"AF",   x"2A",   x"1D",   x"44",   x"73", 
  x"8D",   x"BA",   x"E3",   x"D4",   x"51",   x"66",   x"3F",   x"08", 
  x"2F",   x"18",   x"41",   x"76",   x"F3",   x"C4",   x"9D",   x"AA", 
  x"54",   x"63",   x"3A",   x"0D",   x"88",   x"BF",   x"E6",   x"D1", 
  x"D9",   x"EE",   x"B7",   x"80",   x"05",   x"32",   x"6B",   x"5C", 
  x"A2",   x"95",   x"CC",   x"FB",   x"7E",   x"49",   x"10",   x"27", 
  x"5E",   x"69",   x"30",   x"07",   x"82",   x"B5",   x"EC",   x"DB", 
  x"25",   x"12",   x"4B",   x"7C",   x"F9",   x"CE",   x"97",   x"A0", 
  x"A8",   x"9F",   x"C6",   x"F1",   x"74",   x"43",   x"1A",   x"2D", 
  x"D3",   x"E4",   x"BD",   x"8A",   x"0F",   x"38",   x"61",   x"56", 
  x"71",   x"46",   x"1F",   x"28",   x"AD",   x"9A",   x"C3",   x"F4", 
  x"0A",   x"3D",   x"64",   x"53",   x"D6",   x"E1",   x"B8",   x"8F", 
  x"87",   x"B0",   x"E9",   x"DE",   x"5B",   x"6C",   x"35",   x"02", 
  x"FC",   x"CB",   x"92",   x"A5",   x"20",   x"17",   x"4E",   x"79", 
  x"BC",   x"8B",   x"D2",   x"E5",   x"60",   x"57",   x"0E",   x"39", 
  x"C7",   x"F0",   x"A9",   x"9E",   x"1B",   x"2C",   x"75",   x"42", 
  x"4A",   x"7D",   x"24",   x"13",   x"96",   x"A1",   x"F8",   x"CF", 
  x"31",   x"06",   x"5F",   x"68",   x"ED",   x"DA",   x"83",   x"B4", 
  x"93",   x"A4",   x"FD",   x"CA",   x"4F",   x"78",   x"21",   x"16", 
  x"E8",   x"DF",   x"86",   x"B1",   x"34",   x"03",   x"5A",   x"6D", 
  x"65",   x"52",   x"0B",   x"3C",   x"B9",   x"8E",   x"D7",   x"E0", 
  x"1E",   x"29",   x"70",   x"47",   x"C2",   x"F5",   x"AC",   x"9B", 
  x"E2",   x"D5",   x"8C",   x"BB",   x"3E",   x"09",   x"50",   x"67", 
  x"99",   x"AE",   x"F7",   x"C0",   x"45",   x"72",   x"2B",   x"1C", 
  x"14",   x"23",   x"7A",   x"4D",   x"C8",   x"FF",   x"A6",   x"91", 
  x"6F",   x"58",   x"01",   x"36",   x"B3",   x"84",   x"DD",   x"EA", 
  x"CD",   x"FA",   x"A3",   x"94",   x"11",   x"26",   x"7F",   x"48", 
  x"B6",   x"81",   x"D8",   x"EF",   x"6A",   x"5D",   x"04",   x"33", 
  x"3B",   x"0C",   x"55",   x"62",   x"E7",   x"D0",   x"89",   x"BE", 
  x"40",   x"77",   x"2E",   x"19",   x"9C",   x"AB",   x"F2",   x"C5", 
  x"00",   x"38",   x"70",   x"48",   x"E0",   x"D8",   x"90",   x"A8", 
  x"03",   x"3B",   x"73",   x"4B",   x"E3",   x"DB",   x"93",   x"AB", 
  x"06",   x"3E",   x"76",   x"4E",   x"E6",   x"DE",   x"96",   x"AE", 
  x"05",   x"3D",   x"75",   x"4D",   x"E5",   x"DD",   x"95",   x"AD", 
  x"0C",   x"34",   x"7C",   x"44",   x"EC",   x"D4",   x"9C",   x"A4", 
  x"0F",   x"37",   x"7F",   x"47",   x"EF",   x"D7",   x"9F",   x"A7", 
  x"0A",   x"32",   x"7A",   x"42",   x"EA",   x"D2",   x"9A",   x"A2", 
  x"09",   x"31",   x"79",   x"41",   x"E9",   x"D1",   x"99",   x"A1", 
  x"18",   x"20",   x"68",   x"50",   x"F8",   x"C0",   x"88",   x"B0", 
  x"1B",   x"23",   x"6B",   x"53",   x"FB",   x"C3",   x"8B",   x"B3", 
  x"1E",   x"26",   x"6E",   x"56",   x"FE",   x"C6",   x"8E",   x"B6", 
  x"1D",   x"25",   x"6D",   x"55",   x"FD",   x"C5",   x"8D",   x"B5", 
  x"14",   x"2C",   x"64",   x"5C",   x"F4",   x"CC",   x"84",   x"BC", 
  x"17",   x"2F",   x"67",   x"5F",   x"F7",   x"CF",   x"87",   x"BF", 
  x"12",   x"2A",   x"62",   x"5A",   x"F2",   x"CA",   x"82",   x"BA", 
  x"11",   x"29",   x"61",   x"59",   x"F1",   x"C9",   x"81",   x"B9", 
  x"30",   x"08",   x"40",   x"78",   x"D0",   x"E8",   x"A0",   x"98", 
  x"33",   x"0B",   x"43",   x"7B",   x"D3",   x"EB",   x"A3",   x"9B", 
  x"36",   x"0E",   x"46",   x"7E",   x"D6",   x"EE",   x"A6",   x"9E", 
  x"35",   x"0D",   x"45",   x"7D",   x"D5",   x"ED",   x"A5",   x"9D", 
  x"3C",   x"04",   x"4C",   x"74",   x"DC",   x"E4",   x"AC",   x"94", 
  x"3F",   x"07",   x"4F",   x"77",   x"DF",   x"E7",   x"AF",   x"97", 
  x"3A",   x"02",   x"4A",   x"72",   x"DA",   x"E2",   x"AA",   x"92", 
  x"39",   x"01",   x"49",   x"71",   x"D9",   x"E1",   x"A9",   x"91", 
  x"28",   x"10",   x"58",   x"60",   x"C8",   x"F0",   x"B8",   x"80", 
  x"2B",   x"13",   x"5B",   x"63",   x"CB",   x"F3",   x"BB",   x"83", 
  x"2E",   x"16",   x"5E",   x"66",   x"CE",   x"F6",   x"BE",   x"86", 
  x"2D",   x"15",   x"5D",   x"65",   x"CD",   x"F5",   x"BD",   x"85", 
  x"24",   x"1C",   x"54",   x"6C",   x"C4",   x"FC",   x"B4",   x"8C", 
  x"27",   x"1F",   x"57",   x"6F",   x"C7",   x"FF",   x"B7",   x"8F", 
  x"22",   x"1A",   x"52",   x"6A",   x"C2",   x"FA",   x"B2",   x"8A", 
  x"21",   x"19",   x"51",   x"69",   x"C1",   x"F9",   x"B1",   x"89", 
  x"00",   x"39",   x"72",   x"4B",   x"E4",   x"DD",   x"96",   x"AF", 
  x"0B",   x"32",   x"79",   x"40",   x"EF",   x"D6",   x"9D",   x"A4", 
  x"16",   x"2F",   x"64",   x"5D",   x"F2",   x"CB",   x"80",   x"B9", 
  x"1D",   x"24",   x"6F",   x"56",   x"F9",   x"C0",   x"8B",   x"B2", 
  x"2C",   x"15",   x"5E",   x"67",   x"C8",   x"F1",   x"BA",   x"83", 
  x"27",   x"1E",   x"55",   x"6C",   x"C3",   x"FA",   x"B1",   x"88", 
  x"3A",   x"03",   x"48",   x"71",   x"DE",   x"E7",   x"AC",   x"95", 
  x"31",   x"08",   x"43",   x"7A",   x"D5",   x"EC",   x"A7",   x"9E", 
  x"58",   x"61",   x"2A",   x"13",   x"BC",   x"85",   x"CE",   x"F7", 
  x"53",   x"6A",   x"21",   x"18",   x"B7",   x"8E",   x"C5",   x"FC", 
  x"4E",   x"77",   x"3C",   x"05",   x"AA",   x"93",   x"D8",   x"E1", 
  x"45",   x"7C",   x"37",   x"0E",   x"A1",   x"98",   x"D3",   x"EA", 
  x"74",   x"4D",   x"06",   x"3F",   x"90",   x"A9",   x"E2",   x"DB", 
  x"7F",   x"46",   x"0D",   x"34",   x"9B",   x"A2",   x"E9",   x"D0", 
  x"62",   x"5B",   x"10",   x"29",   x"86",   x"BF",   x"F4",   x"CD", 
  x"69",   x"50",   x"1B",   x"22",   x"8D",   x"B4",   x"FF",   x"C6", 
  x"B0",   x"89",   x"C2",   x"FB",   x"54",   x"6D",   x"26",   x"1F", 
  x"BB",   x"82",   x"C9",   x"F0",   x"5F",   x"66",   x"2D",   x"14", 
  x"A6",   x"9F",   x"D4",   x"ED",   x"42",   x"7B",   x"30",   x"09", 
  x"AD",   x"94",   x"DF",   x"E6",   x"49",   x"70",   x"3B",   x"02", 
  x"9C",   x"A5",   x"EE",   x"D7",   x"78",   x"41",   x"0A",   x"33", 
  x"97",   x"AE",   x"E5",   x"DC",   x"73",   x"4A",   x"01",   x"38", 
  x"8A",   x"B3",   x"F8",   x"C1",   x"6E",   x"57",   x"1C",   x"25", 
  x"81",   x"B8",   x"F3",   x"CA",   x"65",   x"5C",   x"17",   x"2E", 
  x"E8",   x"D1",   x"9A",   x"A3",   x"0C",   x"35",   x"7E",   x"47", 
  x"E3",   x"DA",   x"91",   x"A8",   x"07",   x"3E",   x"75",   x"4C", 
  x"FE",   x"C7",   x"8C",   x"B5",   x"1A",   x"23",   x"68",   x"51", 
  x"F5",   x"CC",   x"87",   x"BE",   x"11",   x"28",   x"63",   x"5A", 
  x"C4",   x"FD",   x"B6",   x"8F",   x"20",   x"19",   x"52",   x"6B", 
  x"CF",   x"F6",   x"BD",   x"84",   x"2B",   x"12",   x"59",   x"60", 
  x"D2",   x"EB",   x"A0",   x"99",   x"36",   x"0F",   x"44",   x"7D", 
  x"D9",   x"E0",   x"AB",   x"92",   x"3D",   x"04",   x"4F",   x"76", 
  x"00",   x"3A",   x"74",   x"4E",   x"E8",   x"D2",   x"9C",   x"A6", 
  x"13",   x"29",   x"67",   x"5D",   x"FB",   x"C1",   x"8F",   x"B5", 
  x"26",   x"1C",   x"52",   x"68",   x"CE",   x"F4",   x"BA",   x"80", 
  x"35",   x"0F",   x"41",   x"7B",   x"DD",   x"E7",   x"A9",   x"93", 
  x"4C",   x"76",   x"38",   x"02",   x"A4",   x"9E",   x"D0",   x"EA", 
  x"5F",   x"65",   x"2B",   x"11",   x"B7",   x"8D",   x"C3",   x"F9", 
  x"6A",   x"50",   x"1E",   x"24",   x"82",   x"B8",   x"F6",   x"CC", 
  x"79",   x"43",   x"0D",   x"37",   x"91",   x"AB",   x"E5",   x"DF", 
  x"98",   x"A2",   x"EC",   x"D6",   x"70",   x"4A",   x"04",   x"3E", 
  x"8B",   x"B1",   x"FF",   x"C5",   x"63",   x"59",   x"17",   x"2D", 
  x"BE",   x"84",   x"CA",   x"F0",   x"56",   x"6C",   x"22",   x"18", 
  x"AD",   x"97",   x"D9",   x"E3",   x"45",   x"7F",   x"31",   x"0B", 
  x"D4",   x"EE",   x"A0",   x"9A",   x"3C",   x"06",   x"48",   x"72", 
  x"C7",   x"FD",   x"B3",   x"89",   x"2F",   x"15",   x"5B",   x"61", 
  x"F2",   x"C8",   x"86",   x"BC",   x"1A",   x"20",   x"6E",   x"54", 
  x"E1",   x"DB",   x"95",   x"AF",   x"09",   x"33",   x"7D",   x"47", 
  x"F3",   x"C9",   x"87",   x"BD",   x"1B",   x"21",   x"6F",   x"55", 
  x"E0",   x"DA",   x"94",   x"AE",   x"08",   x"32",   x"7C",   x"46", 
  x"D5",   x"EF",   x"A1",   x"9B",   x"3D",   x"07",   x"49",   x"73", 
  x"C6",   x"FC",   x"B2",   x"88",   x"2E",   x"14",   x"5A",   x"60", 
  x"BF",   x"85",   x"CB",   x"F1",   x"57",   x"6D",   x"23",   x"19", 
  x"AC",   x"96",   x"D8",   x"E2",   x"44",   x"7E",   x"30",   x"0A", 
  x"99",   x"A3",   x"ED",   x"D7",   x"71",   x"4B",   x"05",   x"3F", 
  x"8A",   x"B0",   x"FE",   x"C4",   x"62",   x"58",   x"16",   x"2C", 
  x"6B",   x"51",   x"1F",   x"25",   x"83",   x"B9",   x"F7",   x"CD", 
  x"78",   x"42",   x"0C",   x"36",   x"90",   x"AA",   x"E4",   x"DE", 
  x"4D",   x"77",   x"39",   x"03",   x"A5",   x"9F",   x"D1",   x"EB", 
  x"5E",   x"64",   x"2A",   x"10",   x"B6",   x"8C",   x"C2",   x"F8", 
  x"27",   x"1D",   x"53",   x"69",   x"CF",   x"F5",   x"BB",   x"81", 
  x"34",   x"0E",   x"40",   x"7A",   x"DC",   x"E6",   x"A8",   x"92", 
  x"01",   x"3B",   x"75",   x"4F",   x"E9",   x"D3",   x"9D",   x"A7", 
  x"12",   x"28",   x"66",   x"5C",   x"FA",   x"C0",   x"8E",   x"B4", 
  x"00",   x"3B",   x"76",   x"4D",   x"EC",   x"D7",   x"9A",   x"A1", 
  x"1B",   x"20",   x"6D",   x"56",   x"F7",   x"CC",   x"81",   x"BA", 
  x"36",   x"0D",   x"40",   x"7B",   x"DA",   x"E1",   x"AC",   x"97", 
  x"2D",   x"16",   x"5B",   x"60",   x"C1",   x"FA",   x"B7",   x"8C", 
  x"6C",   x"57",   x"1A",   x"21",   x"80",   x"BB",   x"F6",   x"CD", 
  x"77",   x"4C",   x"01",   x"3A",   x"9B",   x"A0",   x"ED",   x"D6", 
  x"5A",   x"61",   x"2C",   x"17",   x"B6",   x"8D",   x"C0",   x"FB", 
  x"41",   x"7A",   x"37",   x"0C",   x"AD",   x"96",   x"DB",   x"E0", 
  x"D8",   x"E3",   x"AE",   x"95",   x"34",   x"0F",   x"42",   x"79", 
  x"C3",   x"F8",   x"B5",   x"8E",   x"2F",   x"14",   x"59",   x"62", 
  x"EE",   x"D5",   x"98",   x"A3",   x"02",   x"39",   x"74",   x"4F", 
  x"F5",   x"CE",   x"83",   x"B8",   x"19",   x"22",   x"6F",   x"54", 
  x"B4",   x"8F",   x"C2",   x"F9",   x"58",   x"63",   x"2E",   x"15", 
  x"AF",   x"94",   x"D9",   x"E2",   x"43",   x"78",   x"35",   x"0E", 
  x"82",   x"B9",   x"F4",   x"CF",   x"6E",   x"55",   x"18",   x"23", 
  x"99",   x"A2",   x"EF",   x"D4",   x"75",   x"4E",   x"03",   x"38", 
  x"73",   x"48",   x"05",   x"3E",   x"9F",   x"A4",   x"E9",   x"D2", 
  x"68",   x"53",   x"1E",   x"25",   x"84",   x"BF",   x"F2",   x"C9", 
  x"45",   x"7E",   x"33",   x"08",   x"A9",   x"92",   x"DF",   x"E4", 
  x"5E",   x"65",   x"28",   x"13",   x"B2",   x"89",   x"C4",   x"FF", 
  x"1F",   x"24",   x"69",   x"52",   x"F3",   x"C8",   x"85",   x"BE", 
  x"04",   x"3F",   x"72",   x"49",   x"E8",   x"D3",   x"9E",   x"A5", 
  x"29",   x"12",   x"5F",   x"64",   x"C5",   x"FE",   x"B3",   x"88", 
  x"32",   x"09",   x"44",   x"7F",   x"DE",   x"E5",   x"A8",   x"93", 
  x"AB",   x"90",   x"DD",   x"E6",   x"47",   x"7C",   x"31",   x"0A", 
  x"B0",   x"8B",   x"C6",   x"FD",   x"5C",   x"67",   x"2A",   x"11", 
  x"9D",   x"A6",   x"EB",   x"D0",   x"71",   x"4A",   x"07",   x"3C", 
  x"86",   x"BD",   x"F0",   x"CB",   x"6A",   x"51",   x"1C",   x"27", 
  x"C7",   x"FC",   x"B1",   x"8A",   x"2B",   x"10",   x"5D",   x"66", 
  x"DC",   x"E7",   x"AA",   x"91",   x"30",   x"0B",   x"46",   x"7D", 
  x"F1",   x"CA",   x"87",   x"BC",   x"1D",   x"26",   x"6B",   x"50", 
  x"EA",   x"D1",   x"9C",   x"A7",   x"06",   x"3D",   x"70",   x"4B", 
  x"00",   x"3C",   x"78",   x"44",   x"F0",   x"CC",   x"88",   x"B4", 
  x"23",   x"1F",   x"5B",   x"67",   x"D3",   x"EF",   x"AB",   x"97", 
  x"46",   x"7A",   x"3E",   x"02",   x"B6",   x"8A",   x"CE",   x"F2", 
  x"65",   x"59",   x"1D",   x"21",   x"95",   x"A9",   x"ED",   x"D1", 
  x"8C",   x"B0",   x"F4",   x"C8",   x"7C",   x"40",   x"04",   x"38", 
  x"AF",   x"93",   x"D7",   x"EB",   x"5F",   x"63",   x"27",   x"1B", 
  x"CA",   x"F6",   x"B2",   x"8E",   x"3A",   x"06",   x"42",   x"7E", 
  x"E9",   x"D5",   x"91",   x"AD",   x"19",   x"25",   x"61",   x"5D", 
  x"DB",   x"E7",   x"A3",   x"9F",   x"2B",   x"17",   x"53",   x"6F", 
  x"F8",   x"C4",   x"80",   x"BC",   x"08",   x"34",   x"70",   x"4C", 
  x"9D",   x"A1",   x"E5",   x"D9",   x"6D",   x"51",   x"15",   x"29", 
  x"BE",   x"82",   x"C6",   x"FA",   x"4E",   x"72",   x"36",   x"0A", 
  x"57",   x"6B",   x"2F",   x"13",   x"A7",   x"9B",   x"DF",   x"E3", 
  x"74",   x"48",   x"0C",   x"30",   x"84",   x"B8",   x"FC",   x"C0", 
  x"11",   x"2D",   x"69",   x"55",   x"E1",   x"DD",   x"99",   x"A5", 
  x"32",   x"0E",   x"4A",   x"76",   x"C2",   x"FE",   x"BA",   x"86", 
  x"75",   x"49",   x"0D",   x"31",   x"85",   x"B9",   x"FD",   x"C1", 
  x"56",   x"6A",   x"2E",   x"12",   x"A6",   x"9A",   x"DE",   x"E2", 
  x"33",   x"0F",   x"4B",   x"77",   x"C3",   x"FF",   x"BB",   x"87", 
  x"10",   x"2C",   x"68",   x"54",   x"E0",   x"DC",   x"98",   x"A4", 
  x"F9",   x"C5",   x"81",   x"BD",   x"09",   x"35",   x"71",   x"4D", 
  x"DA",   x"E6",   x"A2",   x"9E",   x"2A",   x"16",   x"52",   x"6E", 
  x"BF",   x"83",   x"C7",   x"FB",   x"4F",   x"73",   x"37",   x"0B", 
  x"9C",   x"A0",   x"E4",   x"D8",   x"6C",   x"50",   x"14",   x"28", 
  x"AE",   x"92",   x"D6",   x"EA",   x"5E",   x"62",   x"26",   x"1A", 
  x"8D",   x"B1",   x"F5",   x"C9",   x"7D",   x"41",   x"05",   x"39", 
  x"E8",   x"D4",   x"90",   x"AC",   x"18",   x"24",   x"60",   x"5C", 
  x"CB",   x"F7",   x"B3",   x"8F",   x"3B",   x"07",   x"43",   x"7F", 
  x"22",   x"1E",   x"5A",   x"66",   x"D2",   x"EE",   x"AA",   x"96", 
  x"01",   x"3D",   x"79",   x"45",   x"F1",   x"CD",   x"89",   x"B5", 
  x"64",   x"58",   x"1C",   x"20",   x"94",   x"A8",   x"EC",   x"D0", 
  x"47",   x"7B",   x"3F",   x"03",   x"B7",   x"8B",   x"CF",   x"F3", 
  x"00",   x"3D",   x"7A",   x"47",   x"F4",   x"C9",   x"8E",   x"B3", 
  x"2B",   x"16",   x"51",   x"6C",   x"DF",   x"E2",   x"A5",   x"98", 
  x"56",   x"6B",   x"2C",   x"11",   x"A2",   x"9F",   x"D8",   x"E5", 
  x"7D",   x"40",   x"07",   x"3A",   x"89",   x"B4",   x"F3",   x"CE", 
  x"AC",   x"91",   x"D6",   x"EB",   x"58",   x"65",   x"22",   x"1F", 
  x"87",   x"BA",   x"FD",   x"C0",   x"73",   x"4E",   x"09",   x"34", 
  x"FA",   x"C7",   x"80",   x"BD",   x"0E",   x"33",   x"74",   x"49", 
  x"D1",   x"EC",   x"AB",   x"96",   x"25",   x"18",   x"5F",   x"62", 
  x"9B",   x"A6",   x"E1",   x"DC",   x"6F",   x"52",   x"15",   x"28", 
  x"B0",   x"8D",   x"CA",   x"F7",   x"44",   x"79",   x"3E",   x"03", 
  x"CD",   x"F0",   x"B7",   x"8A",   x"39",   x"04",   x"43",   x"7E", 
  x"E6",   x"DB",   x"9C",   x"A1",   x"12",   x"2F",   x"68",   x"55", 
  x"37",   x"0A",   x"4D",   x"70",   x"C3",   x"FE",   x"B9",   x"84", 
  x"1C",   x"21",   x"66",   x"5B",   x"E8",   x"D5",   x"92",   x"AF", 
  x"61",   x"5C",   x"1B",   x"26",   x"95",   x"A8",   x"EF",   x"D2", 
  x"4A",   x"77",   x"30",   x"0D",   x"BE",   x"83",   x"C4",   x"F9", 
  x"F5",   x"C8",   x"8F",   x"B2",   x"01",   x"3C",   x"7B",   x"46", 
  x"DE",   x"E3",   x"A4",   x"99",   x"2A",   x"17",   x"50",   x"6D", 
  x"A3",   x"9E",   x"D9",   x"E4",   x"57",   x"6A",   x"2D",   x"10", 
  x"88",   x"B5",   x"F2",   x"CF",   x"7C",   x"41",   x"06",   x"3B", 
  x"59",   x"64",   x"23",   x"1E",   x"AD",   x"90",   x"D7",   x"EA", 
  x"72",   x"4F",   x"08",   x"35",   x"86",   x"BB",   x"FC",   x"C1", 
  x"0F",   x"32",   x"75",   x"48",   x"FB",   x"C6",   x"81",   x"BC", 
  x"24",   x"19",   x"5E",   x"63",   x"D0",   x"ED",   x"AA",   x"97", 
  x"6E",   x"53",   x"14",   x"29",   x"9A",   x"A7",   x"E0",   x"DD", 
  x"45",   x"78",   x"3F",   x"02",   x"B1",   x"8C",   x"CB",   x"F6", 
  x"38",   x"05",   x"42",   x"7F",   x"CC",   x"F1",   x"B6",   x"8B", 
  x"13",   x"2E",   x"69",   x"54",   x"E7",   x"DA",   x"9D",   x"A0", 
  x"C2",   x"FF",   x"B8",   x"85",   x"36",   x"0B",   x"4C",   x"71", 
  x"E9",   x"D4",   x"93",   x"AE",   x"1D",   x"20",   x"67",   x"5A", 
  x"94",   x"A9",   x"EE",   x"D3",   x"60",   x"5D",   x"1A",   x"27", 
  x"BF",   x"82",   x"C5",   x"F8",   x"4B",   x"76",   x"31",   x"0C", 
  x"00",   x"3E",   x"7C",   x"42",   x"F8",   x"C6",   x"84",   x"BA", 
  x"33",   x"0D",   x"4F",   x"71",   x"CB",   x"F5",   x"B7",   x"89", 
  x"66",   x"58",   x"1A",   x"24",   x"9E",   x"A0",   x"E2",   x"DC", 
  x"55",   x"6B",   x"29",   x"17",   x"AD",   x"93",   x"D1",   x"EF", 
  x"CC",   x"F2",   x"B0",   x"8E",   x"34",   x"0A",   x"48",   x"76", 
  x"FF",   x"C1",   x"83",   x"BD",   x"07",   x"39",   x"7B",   x"45", 
  x"AA",   x"94",   x"D6",   x"E8",   x"52",   x"6C",   x"2E",   x"10", 
  x"99",   x"A7",   x"E5",   x"DB",   x"61",   x"5F",   x"1D",   x"23", 
  x"5B",   x"65",   x"27",   x"19",   x"A3",   x"9D",   x"DF",   x"E1", 
  x"68",   x"56",   x"14",   x"2A",   x"90",   x"AE",   x"EC",   x"D2", 
  x"3D",   x"03",   x"41",   x"7F",   x"C5",   x"FB",   x"B9",   x"87", 
  x"0E",   x"30",   x"72",   x"4C",   x"F6",   x"C8",   x"8A",   x"B4", 
  x"97",   x"A9",   x"EB",   x"D5",   x"6F",   x"51",   x"13",   x"2D", 
  x"A4",   x"9A",   x"D8",   x"E6",   x"5C",   x"62",   x"20",   x"1E", 
  x"F1",   x"CF",   x"8D",   x"B3",   x"09",   x"37",   x"75",   x"4B", 
  x"C2",   x"FC",   x"BE",   x"80",   x"3A",   x"04",   x"46",   x"78", 
  x"B6",   x"88",   x"CA",   x"F4",   x"4E",   x"70",   x"32",   x"0C", 
  x"85",   x"BB",   x"F9",   x"C7",   x"7D",   x"43",   x"01",   x"3F", 
  x"D0",   x"EE",   x"AC",   x"92",   x"28",   x"16",   x"54",   x"6A", 
  x"E3",   x"DD",   x"9F",   x"A1",   x"1B",   x"25",   x"67",   x"59", 
  x"7A",   x"44",   x"06",   x"38",   x"82",   x"BC",   x"FE",   x"C0", 
  x"49",   x"77",   x"35",   x"0B",   x"B1",   x"8F",   x"CD",   x"F3", 
  x"1C",   x"22",   x"60",   x"5E",   x"E4",   x"DA",   x"98",   x"A6", 
  x"2F",   x"11",   x"53",   x"6D",   x"D7",   x"E9",   x"AB",   x"95", 
  x"ED",   x"D3",   x"91",   x"AF",   x"15",   x"2B",   x"69",   x"57", 
  x"DE",   x"E0",   x"A2",   x"9C",   x"26",   x"18",   x"5A",   x"64", 
  x"8B",   x"B5",   x"F7",   x"C9",   x"73",   x"4D",   x"0F",   x"31", 
  x"B8",   x"86",   x"C4",   x"FA",   x"40",   x"7E",   x"3C",   x"02", 
  x"21",   x"1F",   x"5D",   x"63",   x"D9",   x"E7",   x"A5",   x"9B", 
  x"12",   x"2C",   x"6E",   x"50",   x"EA",   x"D4",   x"96",   x"A8", 
  x"47",   x"79",   x"3B",   x"05",   x"BF",   x"81",   x"C3",   x"FD", 
  x"74",   x"4A",   x"08",   x"36",   x"8C",   x"B2",   x"F0",   x"CE", 
  x"00",   x"3F",   x"7E",   x"41",   x"FC",   x"C3",   x"82",   x"BD", 
  x"3B",   x"04",   x"45",   x"7A",   x"C7",   x"F8",   x"B9",   x"86", 
  x"76",   x"49",   x"08",   x"37",   x"8A",   x"B5",   x"F4",   x"CB", 
  x"4D",   x"72",   x"33",   x"0C",   x"B1",   x"8E",   x"CF",   x"F0", 
  x"EC",   x"D3",   x"92",   x"AD",   x"10",   x"2F",   x"6E",   x"51", 
  x"D7",   x"E8",   x"A9",   x"96",   x"2B",   x"14",   x"55",   x"6A", 
  x"9A",   x"A5",   x"E4",   x"DB",   x"66",   x"59",   x"18",   x"27", 
  x"A1",   x"9E",   x"DF",   x"E0",   x"5D",   x"62",   x"23",   x"1C", 
  x"1B",   x"24",   x"65",   x"5A",   x"E7",   x"D8",   x"99",   x"A6", 
  x"20",   x"1F",   x"5E",   x"61",   x"DC",   x"E3",   x"A2",   x"9D", 
  x"6D",   x"52",   x"13",   x"2C",   x"91",   x"AE",   x"EF",   x"D0", 
  x"56",   x"69",   x"28",   x"17",   x"AA",   x"95",   x"D4",   x"EB", 
  x"F7",   x"C8",   x"89",   x"B6",   x"0B",   x"34",   x"75",   x"4A", 
  x"CC",   x"F3",   x"B2",   x"8D",   x"30",   x"0F",   x"4E",   x"71", 
  x"81",   x"BE",   x"FF",   x"C0",   x"7D",   x"42",   x"03",   x"3C", 
  x"BA",   x"85",   x"C4",   x"FB",   x"46",   x"79",   x"38",   x"07", 
  x"36",   x"09",   x"48",   x"77",   x"CA",   x"F5",   x"B4",   x"8B", 
  x"0D",   x"32",   x"73",   x"4C",   x"F1",   x"CE",   x"8F",   x"B0", 
  x"40",   x"7F",   x"3E",   x"01",   x"BC",   x"83",   x"C2",   x"FD", 
  x"7B",   x"44",   x"05",   x"3A",   x"87",   x"B8",   x"F9",   x"C6", 
  x"DA",   x"E5",   x"A4",   x"9B",   x"26",   x"19",   x"58",   x"67", 
  x"E1",   x"DE",   x"9F",   x"A0",   x"1D",   x"22",   x"63",   x"5C", 
  x"AC",   x"93",   x"D2",   x"ED",   x"50",   x"6F",   x"2E",   x"11", 
  x"97",   x"A8",   x"E9",   x"D6",   x"6B",   x"54",   x"15",   x"2A", 
  x"2D",   x"12",   x"53",   x"6C",   x"D1",   x"EE",   x"AF",   x"90", 
  x"16",   x"29",   x"68",   x"57",   x"EA",   x"D5",   x"94",   x"AB", 
  x"5B",   x"64",   x"25",   x"1A",   x"A7",   x"98",   x"D9",   x"E6", 
  x"60",   x"5F",   x"1E",   x"21",   x"9C",   x"A3",   x"E2",   x"DD", 
  x"C1",   x"FE",   x"BF",   x"80",   x"3D",   x"02",   x"43",   x"7C", 
  x"FA",   x"C5",   x"84",   x"BB",   x"06",   x"39",   x"78",   x"47", 
  x"B7",   x"88",   x"C9",   x"F6",   x"4B",   x"74",   x"35",   x"0A", 
  x"8C",   x"B3",   x"F2",   x"CD",   x"70",   x"4F",   x"0E",   x"31", 
  x"00",   x"40",   x"80",   x"C0",   x"C3",   x"83",   x"43",   x"03", 
  x"45",   x"05",   x"C5",   x"85",   x"86",   x"C6",   x"06",   x"46", 
  x"8A",   x"CA",   x"0A",   x"4A",   x"49",   x"09",   x"C9",   x"89", 
  x"CF",   x"8F",   x"4F",   x"0F",   x"0C",   x"4C",   x"8C",   x"CC", 
  x"D7",   x"97",   x"57",   x"17",   x"14",   x"54",   x"94",   x"D4", 
  x"92",   x"D2",   x"12",   x"52",   x"51",   x"11",   x"D1",   x"91", 
  x"5D",   x"1D",   x"DD",   x"9D",   x"9E",   x"DE",   x"1E",   x"5E", 
  x"18",   x"58",   x"98",   x"D8",   x"DB",   x"9B",   x"5B",   x"1B", 
  x"6D",   x"2D",   x"ED",   x"AD",   x"AE",   x"EE",   x"2E",   x"6E", 
  x"28",   x"68",   x"A8",   x"E8",   x"EB",   x"AB",   x"6B",   x"2B", 
  x"E7",   x"A7",   x"67",   x"27",   x"24",   x"64",   x"A4",   x"E4", 
  x"A2",   x"E2",   x"22",   x"62",   x"61",   x"21",   x"E1",   x"A1", 
  x"BA",   x"FA",   x"3A",   x"7A",   x"79",   x"39",   x"F9",   x"B9", 
  x"FF",   x"BF",   x"7F",   x"3F",   x"3C",   x"7C",   x"BC",   x"FC", 
  x"30",   x"70",   x"B0",   x"F0",   x"F3",   x"B3",   x"73",   x"33", 
  x"75",   x"35",   x"F5",   x"B5",   x"B6",   x"F6",   x"36",   x"76", 
  x"DA",   x"9A",   x"5A",   x"1A",   x"19",   x"59",   x"99",   x"D9", 
  x"9F",   x"DF",   x"1F",   x"5F",   x"5C",   x"1C",   x"DC",   x"9C", 
  x"50",   x"10",   x"D0",   x"90",   x"93",   x"D3",   x"13",   x"53", 
  x"15",   x"55",   x"95",   x"D5",   x"D6",   x"96",   x"56",   x"16", 
  x"0D",   x"4D",   x"8D",   x"CD",   x"CE",   x"8E",   x"4E",   x"0E", 
  x"48",   x"08",   x"C8",   x"88",   x"8B",   x"CB",   x"0B",   x"4B", 
  x"87",   x"C7",   x"07",   x"47",   x"44",   x"04",   x"C4",   x"84", 
  x"C2",   x"82",   x"42",   x"02",   x"01",   x"41",   x"81",   x"C1", 
  x"B7",   x"F7",   x"37",   x"77",   x"74",   x"34",   x"F4",   x"B4", 
  x"F2",   x"B2",   x"72",   x"32",   x"31",   x"71",   x"B1",   x"F1", 
  x"3D",   x"7D",   x"BD",   x"FD",   x"FE",   x"BE",   x"7E",   x"3E", 
  x"78",   x"38",   x"F8",   x"B8",   x"BB",   x"FB",   x"3B",   x"7B", 
  x"60",   x"20",   x"E0",   x"A0",   x"A3",   x"E3",   x"23",   x"63", 
  x"25",   x"65",   x"A5",   x"E5",   x"E6",   x"A6",   x"66",   x"26", 
  x"EA",   x"AA",   x"6A",   x"2A",   x"29",   x"69",   x"A9",   x"E9", 
  x"AF",   x"EF",   x"2F",   x"6F",   x"6C",   x"2C",   x"EC",   x"AC", 
  x"00",   x"41",   x"82",   x"C3",   x"C7",   x"86",   x"45",   x"04", 
  x"4D",   x"0C",   x"CF",   x"8E",   x"8A",   x"CB",   x"08",   x"49", 
  x"9A",   x"DB",   x"18",   x"59",   x"5D",   x"1C",   x"DF",   x"9E", 
  x"D7",   x"96",   x"55",   x"14",   x"10",   x"51",   x"92",   x"D3", 
  x"F7",   x"B6",   x"75",   x"34",   x"30",   x"71",   x"B2",   x"F3", 
  x"BA",   x"FB",   x"38",   x"79",   x"7D",   x"3C",   x"FF",   x"BE", 
  x"6D",   x"2C",   x"EF",   x"AE",   x"AA",   x"EB",   x"28",   x"69", 
  x"20",   x"61",   x"A2",   x"E3",   x"E7",   x"A6",   x"65",   x"24", 
  x"2D",   x"6C",   x"AF",   x"EE",   x"EA",   x"AB",   x"68",   x"29", 
  x"60",   x"21",   x"E2",   x"A3",   x"A7",   x"E6",   x"25",   x"64", 
  x"B7",   x"F6",   x"35",   x"74",   x"70",   x"31",   x"F2",   x"B3", 
  x"FA",   x"BB",   x"78",   x"39",   x"3D",   x"7C",   x"BF",   x"FE", 
  x"DA",   x"9B",   x"58",   x"19",   x"1D",   x"5C",   x"9F",   x"DE", 
  x"97",   x"D6",   x"15",   x"54",   x"50",   x"11",   x"D2",   x"93", 
  x"40",   x"01",   x"C2",   x"83",   x"87",   x"C6",   x"05",   x"44", 
  x"0D",   x"4C",   x"8F",   x"CE",   x"CA",   x"8B",   x"48",   x"09", 
  x"5A",   x"1B",   x"D8",   x"99",   x"9D",   x"DC",   x"1F",   x"5E", 
  x"17",   x"56",   x"95",   x"D4",   x"D0",   x"91",   x"52",   x"13", 
  x"C0",   x"81",   x"42",   x"03",   x"07",   x"46",   x"85",   x"C4", 
  x"8D",   x"CC",   x"0F",   x"4E",   x"4A",   x"0B",   x"C8",   x"89", 
  x"AD",   x"EC",   x"2F",   x"6E",   x"6A",   x"2B",   x"E8",   x"A9", 
  x"E0",   x"A1",   x"62",   x"23",   x"27",   x"66",   x"A5",   x"E4", 
  x"37",   x"76",   x"B5",   x"F4",   x"F0",   x"B1",   x"72",   x"33", 
  x"7A",   x"3B",   x"F8",   x"B9",   x"BD",   x"FC",   x"3F",   x"7E", 
  x"77",   x"36",   x"F5",   x"B4",   x"B0",   x"F1",   x"32",   x"73", 
  x"3A",   x"7B",   x"B8",   x"F9",   x"FD",   x"BC",   x"7F",   x"3E", 
  x"ED",   x"AC",   x"6F",   x"2E",   x"2A",   x"6B",   x"A8",   x"E9", 
  x"A0",   x"E1",   x"22",   x"63",   x"67",   x"26",   x"E5",   x"A4", 
  x"80",   x"C1",   x"02",   x"43",   x"47",   x"06",   x"C5",   x"84", 
  x"CD",   x"8C",   x"4F",   x"0E",   x"0A",   x"4B",   x"88",   x"C9", 
  x"1A",   x"5B",   x"98",   x"D9",   x"DD",   x"9C",   x"5F",   x"1E", 
  x"57",   x"16",   x"D5",   x"94",   x"90",   x"D1",   x"12",   x"53", 
  x"00",   x"42",   x"84",   x"C6",   x"CB",   x"89",   x"4F",   x"0D", 
  x"55",   x"17",   x"D1",   x"93",   x"9E",   x"DC",   x"1A",   x"58", 
  x"AA",   x"E8",   x"2E",   x"6C",   x"61",   x"23",   x"E5",   x"A7", 
  x"FF",   x"BD",   x"7B",   x"39",   x"34",   x"76",   x"B0",   x"F2", 
  x"97",   x"D5",   x"13",   x"51",   x"5C",   x"1E",   x"D8",   x"9A", 
  x"C2",   x"80",   x"46",   x"04",   x"09",   x"4B",   x"8D",   x"CF", 
  x"3D",   x"7F",   x"B9",   x"FB",   x"F6",   x"B4",   x"72",   x"30", 
  x"68",   x"2A",   x"EC",   x"AE",   x"A3",   x"E1",   x"27",   x"65", 
  x"ED",   x"AF",   x"69",   x"2B",   x"26",   x"64",   x"A2",   x"E0", 
  x"B8",   x"FA",   x"3C",   x"7E",   x"73",   x"31",   x"F7",   x"B5", 
  x"47",   x"05",   x"C3",   x"81",   x"8C",   x"CE",   x"08",   x"4A", 
  x"12",   x"50",   x"96",   x"D4",   x"D9",   x"9B",   x"5D",   x"1F", 
  x"7A",   x"38",   x"FE",   x"BC",   x"B1",   x"F3",   x"35",   x"77", 
  x"2F",   x"6D",   x"AB",   x"E9",   x"E4",   x"A6",   x"60",   x"22", 
  x"D0",   x"92",   x"54",   x"16",   x"1B",   x"59",   x"9F",   x"DD", 
  x"85",   x"C7",   x"01",   x"43",   x"4E",   x"0C",   x"CA",   x"88", 
  x"19",   x"5B",   x"9D",   x"DF",   x"D2",   x"90",   x"56",   x"14", 
  x"4C",   x"0E",   x"C8",   x"8A",   x"87",   x"C5",   x"03",   x"41", 
  x"B3",   x"F1",   x"37",   x"75",   x"78",   x"3A",   x"FC",   x"BE", 
  x"E6",   x"A4",   x"62",   x"20",   x"2D",   x"6F",   x"A9",   x"EB", 
  x"8E",   x"CC",   x"0A",   x"48",   x"45",   x"07",   x"C1",   x"83", 
  x"DB",   x"99",   x"5F",   x"1D",   x"10",   x"52",   x"94",   x"D6", 
  x"24",   x"66",   x"A0",   x"E2",   x"EF",   x"AD",   x"6B",   x"29", 
  x"71",   x"33",   x"F5",   x"B7",   x"BA",   x"F8",   x"3E",   x"7C", 
  x"F4",   x"B6",   x"70",   x"32",   x"3F",   x"7D",   x"BB",   x"F9", 
  x"A1",   x"E3",   x"25",   x"67",   x"6A",   x"28",   x"EE",   x"AC", 
  x"5E",   x"1C",   x"DA",   x"98",   x"95",   x"D7",   x"11",   x"53", 
  x"0B",   x"49",   x"8F",   x"CD",   x"C0",   x"82",   x"44",   x"06", 
  x"63",   x"21",   x"E7",   x"A5",   x"A8",   x"EA",   x"2C",   x"6E", 
  x"36",   x"74",   x"B2",   x"F0",   x"FD",   x"BF",   x"79",   x"3B", 
  x"C9",   x"8B",   x"4D",   x"0F",   x"02",   x"40",   x"86",   x"C4", 
  x"9C",   x"DE",   x"18",   x"5A",   x"57",   x"15",   x"D3",   x"91", 
  x"00",   x"43",   x"86",   x"C5",   x"CF",   x"8C",   x"49",   x"0A", 
  x"5D",   x"1E",   x"DB",   x"98",   x"92",   x"D1",   x"14",   x"57", 
  x"BA",   x"F9",   x"3C",   x"7F",   x"75",   x"36",   x"F3",   x"B0", 
  x"E7",   x"A4",   x"61",   x"22",   x"28",   x"6B",   x"AE",   x"ED", 
  x"B7",   x"F4",   x"31",   x"72",   x"78",   x"3B",   x"FE",   x"BD", 
  x"EA",   x"A9",   x"6C",   x"2F",   x"25",   x"66",   x"A3",   x"E0", 
  x"0D",   x"4E",   x"8B",   x"C8",   x"C2",   x"81",   x"44",   x"07", 
  x"50",   x"13",   x"D6",   x"95",   x"9F",   x"DC",   x"19",   x"5A", 
  x"AD",   x"EE",   x"2B",   x"68",   x"62",   x"21",   x"E4",   x"A7", 
  x"F0",   x"B3",   x"76",   x"35",   x"3F",   x"7C",   x"B9",   x"FA", 
  x"17",   x"54",   x"91",   x"D2",   x"D8",   x"9B",   x"5E",   x"1D", 
  x"4A",   x"09",   x"CC",   x"8F",   x"85",   x"C6",   x"03",   x"40", 
  x"1A",   x"59",   x"9C",   x"DF",   x"D5",   x"96",   x"53",   x"10", 
  x"47",   x"04",   x"C1",   x"82",   x"88",   x"CB",   x"0E",   x"4D", 
  x"A0",   x"E3",   x"26",   x"65",   x"6F",   x"2C",   x"E9",   x"AA", 
  x"FD",   x"BE",   x"7B",   x"38",   x"32",   x"71",   x"B4",   x"F7", 
  x"99",   x"DA",   x"1F",   x"5C",   x"56",   x"15",   x"D0",   x"93", 
  x"C4",   x"87",   x"42",   x"01",   x"0B",   x"48",   x"8D",   x"CE", 
  x"23",   x"60",   x"A5",   x"E6",   x"EC",   x"AF",   x"6A",   x"29", 
  x"7E",   x"3D",   x"F8",   x"BB",   x"B1",   x"F2",   x"37",   x"74", 
  x"2E",   x"6D",   x"A8",   x"EB",   x"E1",   x"A2",   x"67",   x"24", 
  x"73",   x"30",   x"F5",   x"B6",   x"BC",   x"FF",   x"3A",   x"79", 
  x"94",   x"D7",   x"12",   x"51",   x"5B",   x"18",   x"DD",   x"9E", 
  x"C9",   x"8A",   x"4F",   x"0C",   x"06",   x"45",   x"80",   x"C3", 
  x"34",   x"77",   x"B2",   x"F1",   x"FB",   x"B8",   x"7D",   x"3E", 
  x"69",   x"2A",   x"EF",   x"AC",   x"A6",   x"E5",   x"20",   x"63", 
  x"8E",   x"CD",   x"08",   x"4B",   x"41",   x"02",   x"C7",   x"84", 
  x"D3",   x"90",   x"55",   x"16",   x"1C",   x"5F",   x"9A",   x"D9", 
  x"83",   x"C0",   x"05",   x"46",   x"4C",   x"0F",   x"CA",   x"89", 
  x"DE",   x"9D",   x"58",   x"1B",   x"11",   x"52",   x"97",   x"D4", 
  x"39",   x"7A",   x"BF",   x"FC",   x"F6",   x"B5",   x"70",   x"33", 
  x"64",   x"27",   x"E2",   x"A1",   x"AB",   x"E8",   x"2D",   x"6E", 
  x"00",   x"44",   x"88",   x"CC",   x"D3",   x"97",   x"5B",   x"1F", 
  x"65",   x"21",   x"ED",   x"A9",   x"B6",   x"F2",   x"3E",   x"7A", 
  x"CA",   x"8E",   x"42",   x"06",   x"19",   x"5D",   x"91",   x"D5", 
  x"AF",   x"EB",   x"27",   x"63",   x"7C",   x"38",   x"F4",   x"B0", 
  x"57",   x"13",   x"DF",   x"9B",   x"84",   x"C0",   x"0C",   x"48", 
  x"32",   x"76",   x"BA",   x"FE",   x"E1",   x"A5",   x"69",   x"2D", 
  x"9D",   x"D9",   x"15",   x"51",   x"4E",   x"0A",   x"C6",   x"82", 
  x"F8",   x"BC",   x"70",   x"34",   x"2B",   x"6F",   x"A3",   x"E7", 
  x"AE",   x"EA",   x"26",   x"62",   x"7D",   x"39",   x"F5",   x"B1", 
  x"CB",   x"8F",   x"43",   x"07",   x"18",   x"5C",   x"90",   x"D4", 
  x"64",   x"20",   x"EC",   x"A8",   x"B7",   x"F3",   x"3F",   x"7B", 
  x"01",   x"45",   x"89",   x"CD",   x"D2",   x"96",   x"5A",   x"1E", 
  x"F9",   x"BD",   x"71",   x"35",   x"2A",   x"6E",   x"A2",   x"E6", 
  x"9C",   x"D8",   x"14",   x"50",   x"4F",   x"0B",   x"C7",   x"83", 
  x"33",   x"77",   x"BB",   x"FF",   x"E0",   x"A4",   x"68",   x"2C", 
  x"56",   x"12",   x"DE",   x"9A",   x"85",   x"C1",   x"0D",   x"49", 
  x"9F",   x"DB",   x"17",   x"53",   x"4C",   x"08",   x"C4",   x"80", 
  x"FA",   x"BE",   x"72",   x"36",   x"29",   x"6D",   x"A1",   x"E5", 
  x"55",   x"11",   x"DD",   x"99",   x"86",   x"C2",   x"0E",   x"4A", 
  x"30",   x"74",   x"B8",   x"FC",   x"E3",   x"A7",   x"6B",   x"2F", 
  x"C8",   x"8C",   x"40",   x"04",   x"1B",   x"5F",   x"93",   x"D7", 
  x"AD",   x"E9",   x"25",   x"61",   x"7E",   x"3A",   x"F6",   x"B2", 
  x"02",   x"46",   x"8A",   x"CE",   x"D1",   x"95",   x"59",   x"1D", 
  x"67",   x"23",   x"EF",   x"AB",   x"B4",   x"F0",   x"3C",   x"78", 
  x"31",   x"75",   x"B9",   x"FD",   x"E2",   x"A6",   x"6A",   x"2E", 
  x"54",   x"10",   x"DC",   x"98",   x"87",   x"C3",   x"0F",   x"4B", 
  x"FB",   x"BF",   x"73",   x"37",   x"28",   x"6C",   x"A0",   x"E4", 
  x"9E",   x"DA",   x"16",   x"52",   x"4D",   x"09",   x"C5",   x"81", 
  x"66",   x"22",   x"EE",   x"AA",   x"B5",   x"F1",   x"3D",   x"79", 
  x"03",   x"47",   x"8B",   x"CF",   x"D0",   x"94",   x"58",   x"1C", 
  x"AC",   x"E8",   x"24",   x"60",   x"7F",   x"3B",   x"F7",   x"B3", 
  x"C9",   x"8D",   x"41",   x"05",   x"1A",   x"5E",   x"92",   x"D6", 
  x"00",   x"45",   x"8A",   x"CF",   x"D7",   x"92",   x"5D",   x"18", 
  x"6D",   x"28",   x"E7",   x"A2",   x"BA",   x"FF",   x"30",   x"75", 
  x"DA",   x"9F",   x"50",   x"15",   x"0D",   x"48",   x"87",   x"C2", 
  x"B7",   x"F2",   x"3D",   x"78",   x"60",   x"25",   x"EA",   x"AF", 
  x"77",   x"32",   x"FD",   x"B8",   x"A0",   x"E5",   x"2A",   x"6F", 
  x"1A",   x"5F",   x"90",   x"D5",   x"CD",   x"88",   x"47",   x"02", 
  x"AD",   x"E8",   x"27",   x"62",   x"7A",   x"3F",   x"F0",   x"B5", 
  x"C0",   x"85",   x"4A",   x"0F",   x"17",   x"52",   x"9D",   x"D8", 
  x"EE",   x"AB",   x"64",   x"21",   x"39",   x"7C",   x"B3",   x"F6", 
  x"83",   x"C6",   x"09",   x"4C",   x"54",   x"11",   x"DE",   x"9B", 
  x"34",   x"71",   x"BE",   x"FB",   x"E3",   x"A6",   x"69",   x"2C", 
  x"59",   x"1C",   x"D3",   x"96",   x"8E",   x"CB",   x"04",   x"41", 
  x"99",   x"DC",   x"13",   x"56",   x"4E",   x"0B",   x"C4",   x"81", 
  x"F4",   x"B1",   x"7E",   x"3B",   x"23",   x"66",   x"A9",   x"EC", 
  x"43",   x"06",   x"C9",   x"8C",   x"94",   x"D1",   x"1E",   x"5B", 
  x"2E",   x"6B",   x"A4",   x"E1",   x"F9",   x"BC",   x"73",   x"36", 
  x"1F",   x"5A",   x"95",   x"D0",   x"C8",   x"8D",   x"42",   x"07", 
  x"72",   x"37",   x"F8",   x"BD",   x"A5",   x"E0",   x"2F",   x"6A", 
  x"C5",   x"80",   x"4F",   x"0A",   x"12",   x"57",   x"98",   x"DD", 
  x"A8",   x"ED",   x"22",   x"67",   x"7F",   x"3A",   x"F5",   x"B0", 
  x"68",   x"2D",   x"E2",   x"A7",   x"BF",   x"FA",   x"35",   x"70", 
  x"05",   x"40",   x"8F",   x"CA",   x"D2",   x"97",   x"58",   x"1D", 
  x"B2",   x"F7",   x"38",   x"7D",   x"65",   x"20",   x"EF",   x"AA", 
  x"DF",   x"9A",   x"55",   x"10",   x"08",   x"4D",   x"82",   x"C7", 
  x"F1",   x"B4",   x"7B",   x"3E",   x"26",   x"63",   x"AC",   x"E9", 
  x"9C",   x"D9",   x"16",   x"53",   x"4B",   x"0E",   x"C1",   x"84", 
  x"2B",   x"6E",   x"A1",   x"E4",   x"FC",   x"B9",   x"76",   x"33", 
  x"46",   x"03",   x"CC",   x"89",   x"91",   x"D4",   x"1B",   x"5E", 
  x"86",   x"C3",   x"0C",   x"49",   x"51",   x"14",   x"DB",   x"9E", 
  x"EB",   x"AE",   x"61",   x"24",   x"3C",   x"79",   x"B6",   x"F3", 
  x"5C",   x"19",   x"D6",   x"93",   x"8B",   x"CE",   x"01",   x"44", 
  x"31",   x"74",   x"BB",   x"FE",   x"E6",   x"A3",   x"6C",   x"29", 
  x"00",   x"46",   x"8C",   x"CA",   x"DB",   x"9D",   x"57",   x"11", 
  x"75",   x"33",   x"F9",   x"BF",   x"AE",   x"E8",   x"22",   x"64", 
  x"EA",   x"AC",   x"66",   x"20",   x"31",   x"77",   x"BD",   x"FB", 
  x"9F",   x"D9",   x"13",   x"55",   x"44",   x"02",   x"C8",   x"8E", 
  x"17",   x"51",   x"9B",   x"DD",   x"CC",   x"8A",   x"40",   x"06", 
  x"62",   x"24",   x"EE",   x"A8",   x"B9",   x"FF",   x"35",   x"73", 
  x"FD",   x"BB",   x"71",   x"37",   x"26",   x"60",   x"AA",   x"EC", 
  x"88",   x"CE",   x"04",   x"42",   x"53",   x"15",   x"DF",   x"99", 
  x"2E",   x"68",   x"A2",   x"E4",   x"F5",   x"B3",   x"79",   x"3F", 
  x"5B",   x"1D",   x"D7",   x"91",   x"80",   x"C6",   x"0C",   x"4A", 
  x"C4",   x"82",   x"48",   x"0E",   x"1F",   x"59",   x"93",   x"D5", 
  x"B1",   x"F7",   x"3D",   x"7B",   x"6A",   x"2C",   x"E6",   x"A0", 
  x"39",   x"7F",   x"B5",   x"F3",   x"E2",   x"A4",   x"6E",   x"28", 
  x"4C",   x"0A",   x"C0",   x"86",   x"97",   x"D1",   x"1B",   x"5D", 
  x"D3",   x"95",   x"5F",   x"19",   x"08",   x"4E",   x"84",   x"C2", 
  x"A6",   x"E0",   x"2A",   x"6C",   x"7D",   x"3B",   x"F1",   x"B7", 
  x"5C",   x"1A",   x"D0",   x"96",   x"87",   x"C1",   x"0B",   x"4D", 
  x"29",   x"6F",   x"A5",   x"E3",   x"F2",   x"B4",   x"7E",   x"38", 
  x"B6",   x"F0",   x"3A",   x"7C",   x"6D",   x"2B",   x"E1",   x"A7", 
  x"C3",   x"85",   x"4F",   x"09",   x"18",   x"5E",   x"94",   x"D2", 
  x"4B",   x"0D",   x"C7",   x"81",   x"90",   x"D6",   x"1C",   x"5A", 
  x"3E",   x"78",   x"B2",   x"F4",   x"E5",   x"A3",   x"69",   x"2F", 
  x"A1",   x"E7",   x"2D",   x"6B",   x"7A",   x"3C",   x"F6",   x"B0", 
  x"D4",   x"92",   x"58",   x"1E",   x"0F",   x"49",   x"83",   x"C5", 
  x"72",   x"34",   x"FE",   x"B8",   x"A9",   x"EF",   x"25",   x"63", 
  x"07",   x"41",   x"8B",   x"CD",   x"DC",   x"9A",   x"50",   x"16", 
  x"98",   x"DE",   x"14",   x"52",   x"43",   x"05",   x"CF",   x"89", 
  x"ED",   x"AB",   x"61",   x"27",   x"36",   x"70",   x"BA",   x"FC", 
  x"65",   x"23",   x"E9",   x"AF",   x"BE",   x"F8",   x"32",   x"74", 
  x"10",   x"56",   x"9C",   x"DA",   x"CB",   x"8D",   x"47",   x"01", 
  x"8F",   x"C9",   x"03",   x"45",   x"54",   x"12",   x"D8",   x"9E", 
  x"FA",   x"BC",   x"76",   x"30",   x"21",   x"67",   x"AD",   x"EB", 
  x"00",   x"47",   x"8E",   x"C9",   x"DF",   x"98",   x"51",   x"16", 
  x"7D",   x"3A",   x"F3",   x"B4",   x"A2",   x"E5",   x"2C",   x"6B", 
  x"FA",   x"BD",   x"74",   x"33",   x"25",   x"62",   x"AB",   x"EC", 
  x"87",   x"C0",   x"09",   x"4E",   x"58",   x"1F",   x"D6",   x"91", 
  x"37",   x"70",   x"B9",   x"FE",   x"E8",   x"AF",   x"66",   x"21", 
  x"4A",   x"0D",   x"C4",   x"83",   x"95",   x"D2",   x"1B",   x"5C", 
  x"CD",   x"8A",   x"43",   x"04",   x"12",   x"55",   x"9C",   x"DB", 
  x"B0",   x"F7",   x"3E",   x"79",   x"6F",   x"28",   x"E1",   x"A6", 
  x"6E",   x"29",   x"E0",   x"A7",   x"B1",   x"F6",   x"3F",   x"78", 
  x"13",   x"54",   x"9D",   x"DA",   x"CC",   x"8B",   x"42",   x"05", 
  x"94",   x"D3",   x"1A",   x"5D",   x"4B",   x"0C",   x"C5",   x"82", 
  x"E9",   x"AE",   x"67",   x"20",   x"36",   x"71",   x"B8",   x"FF", 
  x"59",   x"1E",   x"D7",   x"90",   x"86",   x"C1",   x"08",   x"4F", 
  x"24",   x"63",   x"AA",   x"ED",   x"FB",   x"BC",   x"75",   x"32", 
  x"A3",   x"E4",   x"2D",   x"6A",   x"7C",   x"3B",   x"F2",   x"B5", 
  x"DE",   x"99",   x"50",   x"17",   x"01",   x"46",   x"8F",   x"C8", 
  x"DC",   x"9B",   x"52",   x"15",   x"03",   x"44",   x"8D",   x"CA", 
  x"A1",   x"E6",   x"2F",   x"68",   x"7E",   x"39",   x"F0",   x"B7", 
  x"26",   x"61",   x"A8",   x"EF",   x"F9",   x"BE",   x"77",   x"30", 
  x"5B",   x"1C",   x"D5",   x"92",   x"84",   x"C3",   x"0A",   x"4D", 
  x"EB",   x"AC",   x"65",   x"22",   x"34",   x"73",   x"BA",   x"FD", 
  x"96",   x"D1",   x"18",   x"5F",   x"49",   x"0E",   x"C7",   x"80", 
  x"11",   x"56",   x"9F",   x"D8",   x"CE",   x"89",   x"40",   x"07", 
  x"6C",   x"2B",   x"E2",   x"A5",   x"B3",   x"F4",   x"3D",   x"7A", 
  x"B2",   x"F5",   x"3C",   x"7B",   x"6D",   x"2A",   x"E3",   x"A4", 
  x"CF",   x"88",   x"41",   x"06",   x"10",   x"57",   x"9E",   x"D9", 
  x"48",   x"0F",   x"C6",   x"81",   x"97",   x"D0",   x"19",   x"5E", 
  x"35",   x"72",   x"BB",   x"FC",   x"EA",   x"AD",   x"64",   x"23", 
  x"85",   x"C2",   x"0B",   x"4C",   x"5A",   x"1D",   x"D4",   x"93", 
  x"F8",   x"BF",   x"76",   x"31",   x"27",   x"60",   x"A9",   x"EE", 
  x"7F",   x"38",   x"F1",   x"B6",   x"A0",   x"E7",   x"2E",   x"69", 
  x"02",   x"45",   x"8C",   x"CB",   x"DD",   x"9A",   x"53",   x"14", 
  x"00",   x"48",   x"90",   x"D8",   x"E3",   x"AB",   x"73",   x"3B", 
  x"05",   x"4D",   x"95",   x"DD",   x"E6",   x"AE",   x"76",   x"3E", 
  x"0A",   x"42",   x"9A",   x"D2",   x"E9",   x"A1",   x"79",   x"31", 
  x"0F",   x"47",   x"9F",   x"D7",   x"EC",   x"A4",   x"7C",   x"34", 
  x"14",   x"5C",   x"84",   x"CC",   x"F7",   x"BF",   x"67",   x"2F", 
  x"11",   x"59",   x"81",   x"C9",   x"F2",   x"BA",   x"62",   x"2A", 
  x"1E",   x"56",   x"8E",   x"C6",   x"FD",   x"B5",   x"6D",   x"25", 
  x"1B",   x"53",   x"8B",   x"C3",   x"F8",   x"B0",   x"68",   x"20", 
  x"28",   x"60",   x"B8",   x"F0",   x"CB",   x"83",   x"5B",   x"13", 
  x"2D",   x"65",   x"BD",   x"F5",   x"CE",   x"86",   x"5E",   x"16", 
  x"22",   x"6A",   x"B2",   x"FA",   x"C1",   x"89",   x"51",   x"19", 
  x"27",   x"6F",   x"B7",   x"FF",   x"C4",   x"8C",   x"54",   x"1C", 
  x"3C",   x"74",   x"AC",   x"E4",   x"DF",   x"97",   x"4F",   x"07", 
  x"39",   x"71",   x"A9",   x"E1",   x"DA",   x"92",   x"4A",   x"02", 
  x"36",   x"7E",   x"A6",   x"EE",   x"D5",   x"9D",   x"45",   x"0D", 
  x"33",   x"7B",   x"A3",   x"EB",   x"D0",   x"98",   x"40",   x"08", 
  x"50",   x"18",   x"C0",   x"88",   x"B3",   x"FB",   x"23",   x"6B", 
  x"55",   x"1D",   x"C5",   x"8D",   x"B6",   x"FE",   x"26",   x"6E", 
  x"5A",   x"12",   x"CA",   x"82",   x"B9",   x"F1",   x"29",   x"61", 
  x"5F",   x"17",   x"CF",   x"87",   x"BC",   x"F4",   x"2C",   x"64", 
  x"44",   x"0C",   x"D4",   x"9C",   x"A7",   x"EF",   x"37",   x"7F", 
  x"41",   x"09",   x"D1",   x"99",   x"A2",   x"EA",   x"32",   x"7A", 
  x"4E",   x"06",   x"DE",   x"96",   x"AD",   x"E5",   x"3D",   x"75", 
  x"4B",   x"03",   x"DB",   x"93",   x"A8",   x"E0",   x"38",   x"70", 
  x"78",   x"30",   x"E8",   x"A0",   x"9B",   x"D3",   x"0B",   x"43", 
  x"7D",   x"35",   x"ED",   x"A5",   x"9E",   x"D6",   x"0E",   x"46", 
  x"72",   x"3A",   x"E2",   x"AA",   x"91",   x"D9",   x"01",   x"49", 
  x"77",   x"3F",   x"E7",   x"AF",   x"94",   x"DC",   x"04",   x"4C", 
  x"6C",   x"24",   x"FC",   x"B4",   x"8F",   x"C7",   x"1F",   x"57", 
  x"69",   x"21",   x"F9",   x"B1",   x"8A",   x"C2",   x"1A",   x"52", 
  x"66",   x"2E",   x"F6",   x"BE",   x"85",   x"CD",   x"15",   x"5D", 
  x"63",   x"2B",   x"F3",   x"BB",   x"80",   x"C8",   x"10",   x"58", 
  x"00",   x"49",   x"92",   x"DB",   x"E7",   x"AE",   x"75",   x"3C", 
  x"0D",   x"44",   x"9F",   x"D6",   x"EA",   x"A3",   x"78",   x"31", 
  x"1A",   x"53",   x"88",   x"C1",   x"FD",   x"B4",   x"6F",   x"26", 
  x"17",   x"5E",   x"85",   x"CC",   x"F0",   x"B9",   x"62",   x"2B", 
  x"34",   x"7D",   x"A6",   x"EF",   x"D3",   x"9A",   x"41",   x"08", 
  x"39",   x"70",   x"AB",   x"E2",   x"DE",   x"97",   x"4C",   x"05", 
  x"2E",   x"67",   x"BC",   x"F5",   x"C9",   x"80",   x"5B",   x"12", 
  x"23",   x"6A",   x"B1",   x"F8",   x"C4",   x"8D",   x"56",   x"1F", 
  x"68",   x"21",   x"FA",   x"B3",   x"8F",   x"C6",   x"1D",   x"54", 
  x"65",   x"2C",   x"F7",   x"BE",   x"82",   x"CB",   x"10",   x"59", 
  x"72",   x"3B",   x"E0",   x"A9",   x"95",   x"DC",   x"07",   x"4E", 
  x"7F",   x"36",   x"ED",   x"A4",   x"98",   x"D1",   x"0A",   x"43", 
  x"5C",   x"15",   x"CE",   x"87",   x"BB",   x"F2",   x"29",   x"60", 
  x"51",   x"18",   x"C3",   x"8A",   x"B6",   x"FF",   x"24",   x"6D", 
  x"46",   x"0F",   x"D4",   x"9D",   x"A1",   x"E8",   x"33",   x"7A", 
  x"4B",   x"02",   x"D9",   x"90",   x"AC",   x"E5",   x"3E",   x"77", 
  x"D0",   x"99",   x"42",   x"0B",   x"37",   x"7E",   x"A5",   x"EC", 
  x"DD",   x"94",   x"4F",   x"06",   x"3A",   x"73",   x"A8",   x"E1", 
  x"CA",   x"83",   x"58",   x"11",   x"2D",   x"64",   x"BF",   x"F6", 
  x"C7",   x"8E",   x"55",   x"1C",   x"20",   x"69",   x"B2",   x"FB", 
  x"E4",   x"AD",   x"76",   x"3F",   x"03",   x"4A",   x"91",   x"D8", 
  x"E9",   x"A0",   x"7B",   x"32",   x"0E",   x"47",   x"9C",   x"D5", 
  x"FE",   x"B7",   x"6C",   x"25",   x"19",   x"50",   x"8B",   x"C2", 
  x"F3",   x"BA",   x"61",   x"28",   x"14",   x"5D",   x"86",   x"CF", 
  x"B8",   x"F1",   x"2A",   x"63",   x"5F",   x"16",   x"CD",   x"84", 
  x"B5",   x"FC",   x"27",   x"6E",   x"52",   x"1B",   x"C0",   x"89", 
  x"A2",   x"EB",   x"30",   x"79",   x"45",   x"0C",   x"D7",   x"9E", 
  x"AF",   x"E6",   x"3D",   x"74",   x"48",   x"01",   x"DA",   x"93", 
  x"8C",   x"C5",   x"1E",   x"57",   x"6B",   x"22",   x"F9",   x"B0", 
  x"81",   x"C8",   x"13",   x"5A",   x"66",   x"2F",   x"F4",   x"BD", 
  x"96",   x"DF",   x"04",   x"4D",   x"71",   x"38",   x"E3",   x"AA", 
  x"9B",   x"D2",   x"09",   x"40",   x"7C",   x"35",   x"EE",   x"A7", 
  x"00",   x"4A",   x"94",   x"DE",   x"EB",   x"A1",   x"7F",   x"35", 
  x"15",   x"5F",   x"81",   x"CB",   x"FE",   x"B4",   x"6A",   x"20", 
  x"2A",   x"60",   x"BE",   x"F4",   x"C1",   x"8B",   x"55",   x"1F", 
  x"3F",   x"75",   x"AB",   x"E1",   x"D4",   x"9E",   x"40",   x"0A", 
  x"54",   x"1E",   x"C0",   x"8A",   x"BF",   x"F5",   x"2B",   x"61", 
  x"41",   x"0B",   x"D5",   x"9F",   x"AA",   x"E0",   x"3E",   x"74", 
  x"7E",   x"34",   x"EA",   x"A0",   x"95",   x"DF",   x"01",   x"4B", 
  x"6B",   x"21",   x"FF",   x"B5",   x"80",   x"CA",   x"14",   x"5E", 
  x"A8",   x"E2",   x"3C",   x"76",   x"43",   x"09",   x"D7",   x"9D", 
  x"BD",   x"F7",   x"29",   x"63",   x"56",   x"1C",   x"C2",   x"88", 
  x"82",   x"C8",   x"16",   x"5C",   x"69",   x"23",   x"FD",   x"B7", 
  x"97",   x"DD",   x"03",   x"49",   x"7C",   x"36",   x"E8",   x"A2", 
  x"FC",   x"B6",   x"68",   x"22",   x"17",   x"5D",   x"83",   x"C9", 
  x"E9",   x"A3",   x"7D",   x"37",   x"02",   x"48",   x"96",   x"DC", 
  x"D6",   x"9C",   x"42",   x"08",   x"3D",   x"77",   x"A9",   x"E3", 
  x"C3",   x"89",   x"57",   x"1D",   x"28",   x"62",   x"BC",   x"F6", 
  x"93",   x"D9",   x"07",   x"4D",   x"78",   x"32",   x"EC",   x"A6", 
  x"86",   x"CC",   x"12",   x"58",   x"6D",   x"27",   x"F9",   x"B3", 
  x"B9",   x"F3",   x"2D",   x"67",   x"52",   x"18",   x"C6",   x"8C", 
  x"AC",   x"E6",   x"38",   x"72",   x"47",   x"0D",   x"D3",   x"99", 
  x"C7",   x"8D",   x"53",   x"19",   x"2C",   x"66",   x"B8",   x"F2", 
  x"D2",   x"98",   x"46",   x"0C",   x"39",   x"73",   x"AD",   x"E7", 
  x"ED",   x"A7",   x"79",   x"33",   x"06",   x"4C",   x"92",   x"D8", 
  x"F8",   x"B2",   x"6C",   x"26",   x"13",   x"59",   x"87",   x"CD", 
  x"3B",   x"71",   x"AF",   x"E5",   x"D0",   x"9A",   x"44",   x"0E", 
  x"2E",   x"64",   x"BA",   x"F0",   x"C5",   x"8F",   x"51",   x"1B", 
  x"11",   x"5B",   x"85",   x"CF",   x"FA",   x"B0",   x"6E",   x"24", 
  x"04",   x"4E",   x"90",   x"DA",   x"EF",   x"A5",   x"7B",   x"31", 
  x"6F",   x"25",   x"FB",   x"B1",   x"84",   x"CE",   x"10",   x"5A", 
  x"7A",   x"30",   x"EE",   x"A4",   x"91",   x"DB",   x"05",   x"4F", 
  x"45",   x"0F",   x"D1",   x"9B",   x"AE",   x"E4",   x"3A",   x"70", 
  x"50",   x"1A",   x"C4",   x"8E",   x"BB",   x"F1",   x"2F",   x"65", 
  x"00",   x"4B",   x"96",   x"DD",   x"EF",   x"A4",   x"79",   x"32", 
  x"1D",   x"56",   x"8B",   x"C0",   x"F2",   x"B9",   x"64",   x"2F", 
  x"3A",   x"71",   x"AC",   x"E7",   x"D5",   x"9E",   x"43",   x"08", 
  x"27",   x"6C",   x"B1",   x"FA",   x"C8",   x"83",   x"5E",   x"15", 
  x"74",   x"3F",   x"E2",   x"A9",   x"9B",   x"D0",   x"0D",   x"46", 
  x"69",   x"22",   x"FF",   x"B4",   x"86",   x"CD",   x"10",   x"5B", 
  x"4E",   x"05",   x"D8",   x"93",   x"A1",   x"EA",   x"37",   x"7C", 
  x"53",   x"18",   x"C5",   x"8E",   x"BC",   x"F7",   x"2A",   x"61", 
  x"E8",   x"A3",   x"7E",   x"35",   x"07",   x"4C",   x"91",   x"DA", 
  x"F5",   x"BE",   x"63",   x"28",   x"1A",   x"51",   x"8C",   x"C7", 
  x"D2",   x"99",   x"44",   x"0F",   x"3D",   x"76",   x"AB",   x"E0", 
  x"CF",   x"84",   x"59",   x"12",   x"20",   x"6B",   x"B6",   x"FD", 
  x"9C",   x"D7",   x"0A",   x"41",   x"73",   x"38",   x"E5",   x"AE", 
  x"81",   x"CA",   x"17",   x"5C",   x"6E",   x"25",   x"F8",   x"B3", 
  x"A6",   x"ED",   x"30",   x"7B",   x"49",   x"02",   x"DF",   x"94", 
  x"BB",   x"F0",   x"2D",   x"66",   x"54",   x"1F",   x"C2",   x"89", 
  x"13",   x"58",   x"85",   x"CE",   x"FC",   x"B7",   x"6A",   x"21", 
  x"0E",   x"45",   x"98",   x"D3",   x"E1",   x"AA",   x"77",   x"3C", 
  x"29",   x"62",   x"BF",   x"F4",   x"C6",   x"8D",   x"50",   x"1B", 
  x"34",   x"7F",   x"A2",   x"E9",   x"DB",   x"90",   x"4D",   x"06", 
  x"67",   x"2C",   x"F1",   x"BA",   x"88",   x"C3",   x"1E",   x"55", 
  x"7A",   x"31",   x"EC",   x"A7",   x"95",   x"DE",   x"03",   x"48", 
  x"5D",   x"16",   x"CB",   x"80",   x"B2",   x"F9",   x"24",   x"6F", 
  x"40",   x"0B",   x"D6",   x"9D",   x"AF",   x"E4",   x"39",   x"72", 
  x"FB",   x"B0",   x"6D",   x"26",   x"14",   x"5F",   x"82",   x"C9", 
  x"E6",   x"AD",   x"70",   x"3B",   x"09",   x"42",   x"9F",   x"D4", 
  x"C1",   x"8A",   x"57",   x"1C",   x"2E",   x"65",   x"B8",   x"F3", 
  x"DC",   x"97",   x"4A",   x"01",   x"33",   x"78",   x"A5",   x"EE", 
  x"8F",   x"C4",   x"19",   x"52",   x"60",   x"2B",   x"F6",   x"BD", 
  x"92",   x"D9",   x"04",   x"4F",   x"7D",   x"36",   x"EB",   x"A0", 
  x"B5",   x"FE",   x"23",   x"68",   x"5A",   x"11",   x"CC",   x"87", 
  x"A8",   x"E3",   x"3E",   x"75",   x"47",   x"0C",   x"D1",   x"9A", 
  x"00",   x"4C",   x"98",   x"D4",   x"F3",   x"BF",   x"6B",   x"27", 
  x"25",   x"69",   x"BD",   x"F1",   x"D6",   x"9A",   x"4E",   x"02", 
  x"4A",   x"06",   x"D2",   x"9E",   x"B9",   x"F5",   x"21",   x"6D", 
  x"6F",   x"23",   x"F7",   x"BB",   x"9C",   x"D0",   x"04",   x"48", 
  x"94",   x"D8",   x"0C",   x"40",   x"67",   x"2B",   x"FF",   x"B3", 
  x"B1",   x"FD",   x"29",   x"65",   x"42",   x"0E",   x"DA",   x"96", 
  x"DE",   x"92",   x"46",   x"0A",   x"2D",   x"61",   x"B5",   x"F9", 
  x"FB",   x"B7",   x"63",   x"2F",   x"08",   x"44",   x"90",   x"DC", 
  x"EB",   x"A7",   x"73",   x"3F",   x"18",   x"54",   x"80",   x"CC", 
  x"CE",   x"82",   x"56",   x"1A",   x"3D",   x"71",   x"A5",   x"E9", 
  x"A1",   x"ED",   x"39",   x"75",   x"52",   x"1E",   x"CA",   x"86", 
  x"84",   x"C8",   x"1C",   x"50",   x"77",   x"3B",   x"EF",   x"A3", 
  x"7F",   x"33",   x"E7",   x"AB",   x"8C",   x"C0",   x"14",   x"58", 
  x"5A",   x"16",   x"C2",   x"8E",   x"A9",   x"E5",   x"31",   x"7D", 
  x"35",   x"79",   x"AD",   x"E1",   x"C6",   x"8A",   x"5E",   x"12", 
  x"10",   x"5C",   x"88",   x"C4",   x"E3",   x"AF",   x"7B",   x"37", 
  x"15",   x"59",   x"8D",   x"C1",   x"E6",   x"AA",   x"7E",   x"32", 
  x"30",   x"7C",   x"A8",   x"E4",   x"C3",   x"8F",   x"5B",   x"17", 
  x"5F",   x"13",   x"C7",   x"8B",   x"AC",   x"E0",   x"34",   x"78", 
  x"7A",   x"36",   x"E2",   x"AE",   x"89",   x"C5",   x"11",   x"5D", 
  x"81",   x"CD",   x"19",   x"55",   x"72",   x"3E",   x"EA",   x"A6", 
  x"A4",   x"E8",   x"3C",   x"70",   x"57",   x"1B",   x"CF",   x"83", 
  x"CB",   x"87",   x"53",   x"1F",   x"38",   x"74",   x"A0",   x"EC", 
  x"EE",   x"A2",   x"76",   x"3A",   x"1D",   x"51",   x"85",   x"C9", 
  x"FE",   x"B2",   x"66",   x"2A",   x"0D",   x"41",   x"95",   x"D9", 
  x"DB",   x"97",   x"43",   x"0F",   x"28",   x"64",   x"B0",   x"FC", 
  x"B4",   x"F8",   x"2C",   x"60",   x"47",   x"0B",   x"DF",   x"93", 
  x"91",   x"DD",   x"09",   x"45",   x"62",   x"2E",   x"FA",   x"B6", 
  x"6A",   x"26",   x"F2",   x"BE",   x"99",   x"D5",   x"01",   x"4D", 
  x"4F",   x"03",   x"D7",   x"9B",   x"BC",   x"F0",   x"24",   x"68", 
  x"20",   x"6C",   x"B8",   x"F4",   x"D3",   x"9F",   x"4B",   x"07", 
  x"05",   x"49",   x"9D",   x"D1",   x"F6",   x"BA",   x"6E",   x"22", 
  x"00",   x"4D",   x"9A",   x"D7",   x"F7",   x"BA",   x"6D",   x"20", 
  x"2D",   x"60",   x"B7",   x"FA",   x"DA",   x"97",   x"40",   x"0D", 
  x"5A",   x"17",   x"C0",   x"8D",   x"AD",   x"E0",   x"37",   x"7A", 
  x"77",   x"3A",   x"ED",   x"A0",   x"80",   x"CD",   x"1A",   x"57", 
  x"B4",   x"F9",   x"2E",   x"63",   x"43",   x"0E",   x"D9",   x"94", 
  x"99",   x"D4",   x"03",   x"4E",   x"6E",   x"23",   x"F4",   x"B9", 
  x"EE",   x"A3",   x"74",   x"39",   x"19",   x"54",   x"83",   x"CE", 
  x"C3",   x"8E",   x"59",   x"14",   x"34",   x"79",   x"AE",   x"E3", 
  x"AB",   x"E6",   x"31",   x"7C",   x"5C",   x"11",   x"C6",   x"8B", 
  x"86",   x"CB",   x"1C",   x"51",   x"71",   x"3C",   x"EB",   x"A6", 
  x"F1",   x"BC",   x"6B",   x"26",   x"06",   x"4B",   x"9C",   x"D1", 
  x"DC",   x"91",   x"46",   x"0B",   x"2B",   x"66",   x"B1",   x"FC", 
  x"1F",   x"52",   x"85",   x"C8",   x"E8",   x"A5",   x"72",   x"3F", 
  x"32",   x"7F",   x"A8",   x"E5",   x"C5",   x"88",   x"5F",   x"12", 
  x"45",   x"08",   x"DF",   x"92",   x"B2",   x"FF",   x"28",   x"65", 
  x"68",   x"25",   x"F2",   x"BF",   x"9F",   x"D2",   x"05",   x"48", 
  x"95",   x"D8",   x"0F",   x"42",   x"62",   x"2F",   x"F8",   x"B5", 
  x"B8",   x"F5",   x"22",   x"6F",   x"4F",   x"02",   x"D5",   x"98", 
  x"CF",   x"82",   x"55",   x"18",   x"38",   x"75",   x"A2",   x"EF", 
  x"E2",   x"AF",   x"78",   x"35",   x"15",   x"58",   x"8F",   x"C2", 
  x"21",   x"6C",   x"BB",   x"F6",   x"D6",   x"9B",   x"4C",   x"01", 
  x"0C",   x"41",   x"96",   x"DB",   x"FB",   x"B6",   x"61",   x"2C", 
  x"7B",   x"36",   x"E1",   x"AC",   x"8C",   x"C1",   x"16",   x"5B", 
  x"56",   x"1B",   x"CC",   x"81",   x"A1",   x"EC",   x"3B",   x"76", 
  x"3E",   x"73",   x"A4",   x"E9",   x"C9",   x"84",   x"53",   x"1E", 
  x"13",   x"5E",   x"89",   x"C4",   x"E4",   x"A9",   x"7E",   x"33", 
  x"64",   x"29",   x"FE",   x"B3",   x"93",   x"DE",   x"09",   x"44", 
  x"49",   x"04",   x"D3",   x"9E",   x"BE",   x"F3",   x"24",   x"69", 
  x"8A",   x"C7",   x"10",   x"5D",   x"7D",   x"30",   x"E7",   x"AA", 
  x"A7",   x"EA",   x"3D",   x"70",   x"50",   x"1D",   x"CA",   x"87", 
  x"D0",   x"9D",   x"4A",   x"07",   x"27",   x"6A",   x"BD",   x"F0", 
  x"FD",   x"B0",   x"67",   x"2A",   x"0A",   x"47",   x"90",   x"DD", 
  x"00",   x"4E",   x"9C",   x"D2",   x"FB",   x"B5",   x"67",   x"29", 
  x"35",   x"7B",   x"A9",   x"E7",   x"CE",   x"80",   x"52",   x"1C", 
  x"6A",   x"24",   x"F6",   x"B8",   x"91",   x"DF",   x"0D",   x"43", 
  x"5F",   x"11",   x"C3",   x"8D",   x"A4",   x"EA",   x"38",   x"76", 
  x"D4",   x"9A",   x"48",   x"06",   x"2F",   x"61",   x"B3",   x"FD", 
  x"E1",   x"AF",   x"7D",   x"33",   x"1A",   x"54",   x"86",   x"C8", 
  x"BE",   x"F0",   x"22",   x"6C",   x"45",   x"0B",   x"D9",   x"97", 
  x"8B",   x"C5",   x"17",   x"59",   x"70",   x"3E",   x"EC",   x"A2", 
  x"6B",   x"25",   x"F7",   x"B9",   x"90",   x"DE",   x"0C",   x"42", 
  x"5E",   x"10",   x"C2",   x"8C",   x"A5",   x"EB",   x"39",   x"77", 
  x"01",   x"4F",   x"9D",   x"D3",   x"FA",   x"B4",   x"66",   x"28", 
  x"34",   x"7A",   x"A8",   x"E6",   x"CF",   x"81",   x"53",   x"1D", 
  x"BF",   x"F1",   x"23",   x"6D",   x"44",   x"0A",   x"D8",   x"96", 
  x"8A",   x"C4",   x"16",   x"58",   x"71",   x"3F",   x"ED",   x"A3", 
  x"D5",   x"9B",   x"49",   x"07",   x"2E",   x"60",   x"B2",   x"FC", 
  x"E0",   x"AE",   x"7C",   x"32",   x"1B",   x"55",   x"87",   x"C9", 
  x"D6",   x"98",   x"4A",   x"04",   x"2D",   x"63",   x"B1",   x"FF", 
  x"E3",   x"AD",   x"7F",   x"31",   x"18",   x"56",   x"84",   x"CA", 
  x"BC",   x"F2",   x"20",   x"6E",   x"47",   x"09",   x"DB",   x"95", 
  x"89",   x"C7",   x"15",   x"5B",   x"72",   x"3C",   x"EE",   x"A0", 
  x"02",   x"4C",   x"9E",   x"D0",   x"F9",   x"B7",   x"65",   x"2B", 
  x"37",   x"79",   x"AB",   x"E5",   x"CC",   x"82",   x"50",   x"1E", 
  x"68",   x"26",   x"F4",   x"BA",   x"93",   x"DD",   x"0F",   x"41", 
  x"5D",   x"13",   x"C1",   x"8F",   x"A6",   x"E8",   x"3A",   x"74", 
  x"BD",   x"F3",   x"21",   x"6F",   x"46",   x"08",   x"DA",   x"94", 
  x"88",   x"C6",   x"14",   x"5A",   x"73",   x"3D",   x"EF",   x"A1", 
  x"D7",   x"99",   x"4B",   x"05",   x"2C",   x"62",   x"B0",   x"FE", 
  x"E2",   x"AC",   x"7E",   x"30",   x"19",   x"57",   x"85",   x"CB", 
  x"69",   x"27",   x"F5",   x"BB",   x"92",   x"DC",   x"0E",   x"40", 
  x"5C",   x"12",   x"C0",   x"8E",   x"A7",   x"E9",   x"3B",   x"75", 
  x"03",   x"4D",   x"9F",   x"D1",   x"F8",   x"B6",   x"64",   x"2A", 
  x"36",   x"78",   x"AA",   x"E4",   x"CD",   x"83",   x"51",   x"1F", 
  x"00",   x"4F",   x"9E",   x"D1",   x"FF",   x"B0",   x"61",   x"2E", 
  x"3D",   x"72",   x"A3",   x"EC",   x"C2",   x"8D",   x"5C",   x"13", 
  x"7A",   x"35",   x"E4",   x"AB",   x"85",   x"CA",   x"1B",   x"54", 
  x"47",   x"08",   x"D9",   x"96",   x"B8",   x"F7",   x"26",   x"69", 
  x"F4",   x"BB",   x"6A",   x"25",   x"0B",   x"44",   x"95",   x"DA", 
  x"C9",   x"86",   x"57",   x"18",   x"36",   x"79",   x"A8",   x"E7", 
  x"8E",   x"C1",   x"10",   x"5F",   x"71",   x"3E",   x"EF",   x"A0", 
  x"B3",   x"FC",   x"2D",   x"62",   x"4C",   x"03",   x"D2",   x"9D", 
  x"2B",   x"64",   x"B5",   x"FA",   x"D4",   x"9B",   x"4A",   x"05", 
  x"16",   x"59",   x"88",   x"C7",   x"E9",   x"A6",   x"77",   x"38", 
  x"51",   x"1E",   x"CF",   x"80",   x"AE",   x"E1",   x"30",   x"7F", 
  x"6C",   x"23",   x"F2",   x"BD",   x"93",   x"DC",   x"0D",   x"42", 
  x"DF",   x"90",   x"41",   x"0E",   x"20",   x"6F",   x"BE",   x"F1", 
  x"E2",   x"AD",   x"7C",   x"33",   x"1D",   x"52",   x"83",   x"CC", 
  x"A5",   x"EA",   x"3B",   x"74",   x"5A",   x"15",   x"C4",   x"8B", 
  x"98",   x"D7",   x"06",   x"49",   x"67",   x"28",   x"F9",   x"B6", 
  x"56",   x"19",   x"C8",   x"87",   x"A9",   x"E6",   x"37",   x"78", 
  x"6B",   x"24",   x"F5",   x"BA",   x"94",   x"DB",   x"0A",   x"45", 
  x"2C",   x"63",   x"B2",   x"FD",   x"D3",   x"9C",   x"4D",   x"02", 
  x"11",   x"5E",   x"8F",   x"C0",   x"EE",   x"A1",   x"70",   x"3F", 
  x"A2",   x"ED",   x"3C",   x"73",   x"5D",   x"12",   x"C3",   x"8C", 
  x"9F",   x"D0",   x"01",   x"4E",   x"60",   x"2F",   x"FE",   x"B1", 
  x"D8",   x"97",   x"46",   x"09",   x"27",   x"68",   x"B9",   x"F6", 
  x"E5",   x"AA",   x"7B",   x"34",   x"1A",   x"55",   x"84",   x"CB", 
  x"7D",   x"32",   x"E3",   x"AC",   x"82",   x"CD",   x"1C",   x"53", 
  x"40",   x"0F",   x"DE",   x"91",   x"BF",   x"F0",   x"21",   x"6E", 
  x"07",   x"48",   x"99",   x"D6",   x"F8",   x"B7",   x"66",   x"29", 
  x"3A",   x"75",   x"A4",   x"EB",   x"C5",   x"8A",   x"5B",   x"14", 
  x"89",   x"C6",   x"17",   x"58",   x"76",   x"39",   x"E8",   x"A7", 
  x"B4",   x"FB",   x"2A",   x"65",   x"4B",   x"04",   x"D5",   x"9A", 
  x"F3",   x"BC",   x"6D",   x"22",   x"0C",   x"43",   x"92",   x"DD", 
  x"CE",   x"81",   x"50",   x"1F",   x"31",   x"7E",   x"AF",   x"E0", 
  x"00",   x"50",   x"A0",   x"F0",   x"83",   x"D3",   x"23",   x"73", 
  x"C5",   x"95",   x"65",   x"35",   x"46",   x"16",   x"E6",   x"B6", 
  x"49",   x"19",   x"E9",   x"B9",   x"CA",   x"9A",   x"6A",   x"3A", 
  x"8C",   x"DC",   x"2C",   x"7C",   x"0F",   x"5F",   x"AF",   x"FF", 
  x"92",   x"C2",   x"32",   x"62",   x"11",   x"41",   x"B1",   x"E1", 
  x"57",   x"07",   x"F7",   x"A7",   x"D4",   x"84",   x"74",   x"24", 
  x"DB",   x"8B",   x"7B",   x"2B",   x"58",   x"08",   x"F8",   x"A8", 
  x"1E",   x"4E",   x"BE",   x"EE",   x"9D",   x"CD",   x"3D",   x"6D", 
  x"E7",   x"B7",   x"47",   x"17",   x"64",   x"34",   x"C4",   x"94", 
  x"22",   x"72",   x"82",   x"D2",   x"A1",   x"F1",   x"01",   x"51", 
  x"AE",   x"FE",   x"0E",   x"5E",   x"2D",   x"7D",   x"8D",   x"DD", 
  x"6B",   x"3B",   x"CB",   x"9B",   x"E8",   x"B8",   x"48",   x"18", 
  x"75",   x"25",   x"D5",   x"85",   x"F6",   x"A6",   x"56",   x"06", 
  x"B0",   x"E0",   x"10",   x"40",   x"33",   x"63",   x"93",   x"C3", 
  x"3C",   x"6C",   x"9C",   x"CC",   x"BF",   x"EF",   x"1F",   x"4F", 
  x"F9",   x"A9",   x"59",   x"09",   x"7A",   x"2A",   x"DA",   x"8A", 
  x"0D",   x"5D",   x"AD",   x"FD",   x"8E",   x"DE",   x"2E",   x"7E", 
  x"C8",   x"98",   x"68",   x"38",   x"4B",   x"1B",   x"EB",   x"BB", 
  x"44",   x"14",   x"E4",   x"B4",   x"C7",   x"97",   x"67",   x"37", 
  x"81",   x"D1",   x"21",   x"71",   x"02",   x"52",   x"A2",   x"F2", 
  x"9F",   x"CF",   x"3F",   x"6F",   x"1C",   x"4C",   x"BC",   x"EC", 
  x"5A",   x"0A",   x"FA",   x"AA",   x"D9",   x"89",   x"79",   x"29", 
  x"D6",   x"86",   x"76",   x"26",   x"55",   x"05",   x"F5",   x"A5", 
  x"13",   x"43",   x"B3",   x"E3",   x"90",   x"C0",   x"30",   x"60", 
  x"EA",   x"BA",   x"4A",   x"1A",   x"69",   x"39",   x"C9",   x"99", 
  x"2F",   x"7F",   x"8F",   x"DF",   x"AC",   x"FC",   x"0C",   x"5C", 
  x"A3",   x"F3",   x"03",   x"53",   x"20",   x"70",   x"80",   x"D0", 
  x"66",   x"36",   x"C6",   x"96",   x"E5",   x"B5",   x"45",   x"15", 
  x"78",   x"28",   x"D8",   x"88",   x"FB",   x"AB",   x"5B",   x"0B", 
  x"BD",   x"ED",   x"1D",   x"4D",   x"3E",   x"6E",   x"9E",   x"CE", 
  x"31",   x"61",   x"91",   x"C1",   x"B2",   x"E2",   x"12",   x"42", 
  x"F4",   x"A4",   x"54",   x"04",   x"77",   x"27",   x"D7",   x"87", 
  x"00",   x"51",   x"A2",   x"F3",   x"87",   x"D6",   x"25",   x"74", 
  x"CD",   x"9C",   x"6F",   x"3E",   x"4A",   x"1B",   x"E8",   x"B9", 
  x"59",   x"08",   x"FB",   x"AA",   x"DE",   x"8F",   x"7C",   x"2D", 
  x"94",   x"C5",   x"36",   x"67",   x"13",   x"42",   x"B1",   x"E0", 
  x"B2",   x"E3",   x"10",   x"41",   x"35",   x"64",   x"97",   x"C6", 
  x"7F",   x"2E",   x"DD",   x"8C",   x"F8",   x"A9",   x"5A",   x"0B", 
  x"EB",   x"BA",   x"49",   x"18",   x"6C",   x"3D",   x"CE",   x"9F", 
  x"26",   x"77",   x"84",   x"D5",   x"A1",   x"F0",   x"03",   x"52", 
  x"A7",   x"F6",   x"05",   x"54",   x"20",   x"71",   x"82",   x"D3", 
  x"6A",   x"3B",   x"C8",   x"99",   x"ED",   x"BC",   x"4F",   x"1E", 
  x"FE",   x"AF",   x"5C",   x"0D",   x"79",   x"28",   x"DB",   x"8A", 
  x"33",   x"62",   x"91",   x"C0",   x"B4",   x"E5",   x"16",   x"47", 
  x"15",   x"44",   x"B7",   x"E6",   x"92",   x"C3",   x"30",   x"61", 
  x"D8",   x"89",   x"7A",   x"2B",   x"5F",   x"0E",   x"FD",   x"AC", 
  x"4C",   x"1D",   x"EE",   x"BF",   x"CB",   x"9A",   x"69",   x"38", 
  x"81",   x"D0",   x"23",   x"72",   x"06",   x"57",   x"A4",   x"F5", 
  x"8D",   x"DC",   x"2F",   x"7E",   x"0A",   x"5B",   x"A8",   x"F9", 
  x"40",   x"11",   x"E2",   x"B3",   x"C7",   x"96",   x"65",   x"34", 
  x"D4",   x"85",   x"76",   x"27",   x"53",   x"02",   x"F1",   x"A0", 
  x"19",   x"48",   x"BB",   x"EA",   x"9E",   x"CF",   x"3C",   x"6D", 
  x"3F",   x"6E",   x"9D",   x"CC",   x"B8",   x"E9",   x"1A",   x"4B", 
  x"F2",   x"A3",   x"50",   x"01",   x"75",   x"24",   x"D7",   x"86", 
  x"66",   x"37",   x"C4",   x"95",   x"E1",   x"B0",   x"43",   x"12", 
  x"AB",   x"FA",   x"09",   x"58",   x"2C",   x"7D",   x"8E",   x"DF", 
  x"2A",   x"7B",   x"88",   x"D9",   x"AD",   x"FC",   x"0F",   x"5E", 
  x"E7",   x"B6",   x"45",   x"14",   x"60",   x"31",   x"C2",   x"93", 
  x"73",   x"22",   x"D1",   x"80",   x"F4",   x"A5",   x"56",   x"07", 
  x"BE",   x"EF",   x"1C",   x"4D",   x"39",   x"68",   x"9B",   x"CA", 
  x"98",   x"C9",   x"3A",   x"6B",   x"1F",   x"4E",   x"BD",   x"EC", 
  x"55",   x"04",   x"F7",   x"A6",   x"D2",   x"83",   x"70",   x"21", 
  x"C1",   x"90",   x"63",   x"32",   x"46",   x"17",   x"E4",   x"B5", 
  x"0C",   x"5D",   x"AE",   x"FF",   x"8B",   x"DA",   x"29",   x"78", 
  x"00",   x"52",   x"A4",   x"F6",   x"8B",   x"D9",   x"2F",   x"7D", 
  x"D5",   x"87",   x"71",   x"23",   x"5E",   x"0C",   x"FA",   x"A8", 
  x"69",   x"3B",   x"CD",   x"9F",   x"E2",   x"B0",   x"46",   x"14", 
  x"BC",   x"EE",   x"18",   x"4A",   x"37",   x"65",   x"93",   x"C1", 
  x"D2",   x"80",   x"76",   x"24",   x"59",   x"0B",   x"FD",   x"AF", 
  x"07",   x"55",   x"A3",   x"F1",   x"8C",   x"DE",   x"28",   x"7A", 
  x"BB",   x"E9",   x"1F",   x"4D",   x"30",   x"62",   x"94",   x"C6", 
  x"6E",   x"3C",   x"CA",   x"98",   x"E5",   x"B7",   x"41",   x"13", 
  x"67",   x"35",   x"C3",   x"91",   x"EC",   x"BE",   x"48",   x"1A", 
  x"B2",   x"E0",   x"16",   x"44",   x"39",   x"6B",   x"9D",   x"CF", 
  x"0E",   x"5C",   x"AA",   x"F8",   x"85",   x"D7",   x"21",   x"73", 
  x"DB",   x"89",   x"7F",   x"2D",   x"50",   x"02",   x"F4",   x"A6", 
  x"B5",   x"E7",   x"11",   x"43",   x"3E",   x"6C",   x"9A",   x"C8", 
  x"60",   x"32",   x"C4",   x"96",   x"EB",   x"B9",   x"4F",   x"1D", 
  x"DC",   x"8E",   x"78",   x"2A",   x"57",   x"05",   x"F3",   x"A1", 
  x"09",   x"5B",   x"AD",   x"FF",   x"82",   x"D0",   x"26",   x"74", 
  x"CE",   x"9C",   x"6A",   x"38",   x"45",   x"17",   x"E1",   x"B3", 
  x"1B",   x"49",   x"BF",   x"ED",   x"90",   x"C2",   x"34",   x"66", 
  x"A7",   x"F5",   x"03",   x"51",   x"2C",   x"7E",   x"88",   x"DA", 
  x"72",   x"20",   x"D6",   x"84",   x"F9",   x"AB",   x"5D",   x"0F", 
  x"1C",   x"4E",   x"B8",   x"EA",   x"97",   x"C5",   x"33",   x"61", 
  x"C9",   x"9B",   x"6D",   x"3F",   x"42",   x"10",   x"E6",   x"B4", 
  x"75",   x"27",   x"D1",   x"83",   x"FE",   x"AC",   x"5A",   x"08", 
  x"A0",   x"F2",   x"04",   x"56",   x"2B",   x"79",   x"8F",   x"DD", 
  x"A9",   x"FB",   x"0D",   x"5F",   x"22",   x"70",   x"86",   x"D4", 
  x"7C",   x"2E",   x"D8",   x"8A",   x"F7",   x"A5",   x"53",   x"01", 
  x"C0",   x"92",   x"64",   x"36",   x"4B",   x"19",   x"EF",   x"BD", 
  x"15",   x"47",   x"B1",   x"E3",   x"9E",   x"CC",   x"3A",   x"68", 
  x"7B",   x"29",   x"DF",   x"8D",   x"F0",   x"A2",   x"54",   x"06", 
  x"AE",   x"FC",   x"0A",   x"58",   x"25",   x"77",   x"81",   x"D3", 
  x"12",   x"40",   x"B6",   x"E4",   x"99",   x"CB",   x"3D",   x"6F", 
  x"C7",   x"95",   x"63",   x"31",   x"4C",   x"1E",   x"E8",   x"BA", 
  x"00",   x"53",   x"A6",   x"F5",   x"8F",   x"DC",   x"29",   x"7A", 
  x"DD",   x"8E",   x"7B",   x"28",   x"52",   x"01",   x"F4",   x"A7", 
  x"79",   x"2A",   x"DF",   x"8C",   x"F6",   x"A5",   x"50",   x"03", 
  x"A4",   x"F7",   x"02",   x"51",   x"2B",   x"78",   x"8D",   x"DE", 
  x"F2",   x"A1",   x"54",   x"07",   x"7D",   x"2E",   x"DB",   x"88", 
  x"2F",   x"7C",   x"89",   x"DA",   x"A0",   x"F3",   x"06",   x"55", 
  x"8B",   x"D8",   x"2D",   x"7E",   x"04",   x"57",   x"A2",   x"F1", 
  x"56",   x"05",   x"F0",   x"A3",   x"D9",   x"8A",   x"7F",   x"2C", 
  x"27",   x"74",   x"81",   x"D2",   x"A8",   x"FB",   x"0E",   x"5D", 
  x"FA",   x"A9",   x"5C",   x"0F",   x"75",   x"26",   x"D3",   x"80", 
  x"5E",   x"0D",   x"F8",   x"AB",   x"D1",   x"82",   x"77",   x"24", 
  x"83",   x"D0",   x"25",   x"76",   x"0C",   x"5F",   x"AA",   x"F9", 
  x"D5",   x"86",   x"73",   x"20",   x"5A",   x"09",   x"FC",   x"AF", 
  x"08",   x"5B",   x"AE",   x"FD",   x"87",   x"D4",   x"21",   x"72", 
  x"AC",   x"FF",   x"0A",   x"59",   x"23",   x"70",   x"85",   x"D6", 
  x"71",   x"22",   x"D7",   x"84",   x"FE",   x"AD",   x"58",   x"0B", 
  x"4E",   x"1D",   x"E8",   x"BB",   x"C1",   x"92",   x"67",   x"34", 
  x"93",   x"C0",   x"35",   x"66",   x"1C",   x"4F",   x"BA",   x"E9", 
  x"37",   x"64",   x"91",   x"C2",   x"B8",   x"EB",   x"1E",   x"4D", 
  x"EA",   x"B9",   x"4C",   x"1F",   x"65",   x"36",   x"C3",   x"90", 
  x"BC",   x"EF",   x"1A",   x"49",   x"33",   x"60",   x"95",   x"C6", 
  x"61",   x"32",   x"C7",   x"94",   x"EE",   x"BD",   x"48",   x"1B", 
  x"C5",   x"96",   x"63",   x"30",   x"4A",   x"19",   x"EC",   x"BF", 
  x"18",   x"4B",   x"BE",   x"ED",   x"97",   x"C4",   x"31",   x"62", 
  x"69",   x"3A",   x"CF",   x"9C",   x"E6",   x"B5",   x"40",   x"13", 
  x"B4",   x"E7",   x"12",   x"41",   x"3B",   x"68",   x"9D",   x"CE", 
  x"10",   x"43",   x"B6",   x"E5",   x"9F",   x"CC",   x"39",   x"6A", 
  x"CD",   x"9E",   x"6B",   x"38",   x"42",   x"11",   x"E4",   x"B7", 
  x"9B",   x"C8",   x"3D",   x"6E",   x"14",   x"47",   x"B2",   x"E1", 
  x"46",   x"15",   x"E0",   x"B3",   x"C9",   x"9A",   x"6F",   x"3C", 
  x"E2",   x"B1",   x"44",   x"17",   x"6D",   x"3E",   x"CB",   x"98", 
  x"3F",   x"6C",   x"99",   x"CA",   x"B0",   x"E3",   x"16",   x"45", 
  x"00",   x"54",   x"A8",   x"FC",   x"93",   x"C7",   x"3B",   x"6F", 
  x"E5",   x"B1",   x"4D",   x"19",   x"76",   x"22",   x"DE",   x"8A", 
  x"09",   x"5D",   x"A1",   x"F5",   x"9A",   x"CE",   x"32",   x"66", 
  x"EC",   x"B8",   x"44",   x"10",   x"7F",   x"2B",   x"D7",   x"83", 
  x"12",   x"46",   x"BA",   x"EE",   x"81",   x"D5",   x"29",   x"7D", 
  x"F7",   x"A3",   x"5F",   x"0B",   x"64",   x"30",   x"CC",   x"98", 
  x"1B",   x"4F",   x"B3",   x"E7",   x"88",   x"DC",   x"20",   x"74", 
  x"FE",   x"AA",   x"56",   x"02",   x"6D",   x"39",   x"C5",   x"91", 
  x"24",   x"70",   x"8C",   x"D8",   x"B7",   x"E3",   x"1F",   x"4B", 
  x"C1",   x"95",   x"69",   x"3D",   x"52",   x"06",   x"FA",   x"AE", 
  x"2D",   x"79",   x"85",   x"D1",   x"BE",   x"EA",   x"16",   x"42", 
  x"C8",   x"9C",   x"60",   x"34",   x"5B",   x"0F",   x"F3",   x"A7", 
  x"36",   x"62",   x"9E",   x"CA",   x"A5",   x"F1",   x"0D",   x"59", 
  x"D3",   x"87",   x"7B",   x"2F",   x"40",   x"14",   x"E8",   x"BC", 
  x"3F",   x"6B",   x"97",   x"C3",   x"AC",   x"F8",   x"04",   x"50", 
  x"DA",   x"8E",   x"72",   x"26",   x"49",   x"1D",   x"E1",   x"B5", 
  x"48",   x"1C",   x"E0",   x"B4",   x"DB",   x"8F",   x"73",   x"27", 
  x"AD",   x"F9",   x"05",   x"51",   x"3E",   x"6A",   x"96",   x"C2", 
  x"41",   x"15",   x"E9",   x"BD",   x"D2",   x"86",   x"7A",   x"2E", 
  x"A4",   x"F0",   x"0C",   x"58",   x"37",   x"63",   x"9F",   x"CB", 
  x"5A",   x"0E",   x"F2",   x"A6",   x"C9",   x"9D",   x"61",   x"35", 
  x"BF",   x"EB",   x"17",   x"43",   x"2C",   x"78",   x"84",   x"D0", 
  x"53",   x"07",   x"FB",   x"AF",   x"C0",   x"94",   x"68",   x"3C", 
  x"B6",   x"E2",   x"1E",   x"4A",   x"25",   x"71",   x"8D",   x"D9", 
  x"6C",   x"38",   x"C4",   x"90",   x"FF",   x"AB",   x"57",   x"03", 
  x"89",   x"DD",   x"21",   x"75",   x"1A",   x"4E",   x"B2",   x"E6", 
  x"65",   x"31",   x"CD",   x"99",   x"F6",   x"A2",   x"5E",   x"0A", 
  x"80",   x"D4",   x"28",   x"7C",   x"13",   x"47",   x"BB",   x"EF", 
  x"7E",   x"2A",   x"D6",   x"82",   x"ED",   x"B9",   x"45",   x"11", 
  x"9B",   x"CF",   x"33",   x"67",   x"08",   x"5C",   x"A0",   x"F4", 
  x"77",   x"23",   x"DF",   x"8B",   x"E4",   x"B0",   x"4C",   x"18", 
  x"92",   x"C6",   x"3A",   x"6E",   x"01",   x"55",   x"A9",   x"FD", 
  x"00",   x"55",   x"AA",   x"FF",   x"97",   x"C2",   x"3D",   x"68", 
  x"ED",   x"B8",   x"47",   x"12",   x"7A",   x"2F",   x"D0",   x"85", 
  x"19",   x"4C",   x"B3",   x"E6",   x"8E",   x"DB",   x"24",   x"71", 
  x"F4",   x"A1",   x"5E",   x"0B",   x"63",   x"36",   x"C9",   x"9C", 
  x"32",   x"67",   x"98",   x"CD",   x"A5",   x"F0",   x"0F",   x"5A", 
  x"DF",   x"8A",   x"75",   x"20",   x"48",   x"1D",   x"E2",   x"B7", 
  x"2B",   x"7E",   x"81",   x"D4",   x"BC",   x"E9",   x"16",   x"43", 
  x"C6",   x"93",   x"6C",   x"39",   x"51",   x"04",   x"FB",   x"AE", 
  x"64",   x"31",   x"CE",   x"9B",   x"F3",   x"A6",   x"59",   x"0C", 
  x"89",   x"DC",   x"23",   x"76",   x"1E",   x"4B",   x"B4",   x"E1", 
  x"7D",   x"28",   x"D7",   x"82",   x"EA",   x"BF",   x"40",   x"15", 
  x"90",   x"C5",   x"3A",   x"6F",   x"07",   x"52",   x"AD",   x"F8", 
  x"56",   x"03",   x"FC",   x"A9",   x"C1",   x"94",   x"6B",   x"3E", 
  x"BB",   x"EE",   x"11",   x"44",   x"2C",   x"79",   x"86",   x"D3", 
  x"4F",   x"1A",   x"E5",   x"B0",   x"D8",   x"8D",   x"72",   x"27", 
  x"A2",   x"F7",   x"08",   x"5D",   x"35",   x"60",   x"9F",   x"CA", 
  x"C8",   x"9D",   x"62",   x"37",   x"5F",   x"0A",   x"F5",   x"A0", 
  x"25",   x"70",   x"8F",   x"DA",   x"B2",   x"E7",   x"18",   x"4D", 
  x"D1",   x"84",   x"7B",   x"2E",   x"46",   x"13",   x"EC",   x"B9", 
  x"3C",   x"69",   x"96",   x"C3",   x"AB",   x"FE",   x"01",   x"54", 
  x"FA",   x"AF",   x"50",   x"05",   x"6D",   x"38",   x"C7",   x"92", 
  x"17",   x"42",   x"BD",   x"E8",   x"80",   x"D5",   x"2A",   x"7F", 
  x"E3",   x"B6",   x"49",   x"1C",   x"74",   x"21",   x"DE",   x"8B", 
  x"0E",   x"5B",   x"A4",   x"F1",   x"99",   x"CC",   x"33",   x"66", 
  x"AC",   x"F9",   x"06",   x"53",   x"3B",   x"6E",   x"91",   x"C4", 
  x"41",   x"14",   x"EB",   x"BE",   x"D6",   x"83",   x"7C",   x"29", 
  x"B5",   x"E0",   x"1F",   x"4A",   x"22",   x"77",   x"88",   x"DD", 
  x"58",   x"0D",   x"F2",   x"A7",   x"CF",   x"9A",   x"65",   x"30", 
  x"9E",   x"CB",   x"34",   x"61",   x"09",   x"5C",   x"A3",   x"F6", 
  x"73",   x"26",   x"D9",   x"8C",   x"E4",   x"B1",   x"4E",   x"1B", 
  x"87",   x"D2",   x"2D",   x"78",   x"10",   x"45",   x"BA",   x"EF", 
  x"6A",   x"3F",   x"C0",   x"95",   x"FD",   x"A8",   x"57",   x"02", 
  x"00",   x"56",   x"AC",   x"FA",   x"9B",   x"CD",   x"37",   x"61", 
  x"F5",   x"A3",   x"59",   x"0F",   x"6E",   x"38",   x"C2",   x"94", 
  x"29",   x"7F",   x"85",   x"D3",   x"B2",   x"E4",   x"1E",   x"48", 
  x"DC",   x"8A",   x"70",   x"26",   x"47",   x"11",   x"EB",   x"BD", 
  x"52",   x"04",   x"FE",   x"A8",   x"C9",   x"9F",   x"65",   x"33", 
  x"A7",   x"F1",   x"0B",   x"5D",   x"3C",   x"6A",   x"90",   x"C6", 
  x"7B",   x"2D",   x"D7",   x"81",   x"E0",   x"B6",   x"4C",   x"1A", 
  x"8E",   x"D8",   x"22",   x"74",   x"15",   x"43",   x"B9",   x"EF", 
  x"A4",   x"F2",   x"08",   x"5E",   x"3F",   x"69",   x"93",   x"C5", 
  x"51",   x"07",   x"FD",   x"AB",   x"CA",   x"9C",   x"66",   x"30", 
  x"8D",   x"DB",   x"21",   x"77",   x"16",   x"40",   x"BA",   x"EC", 
  x"78",   x"2E",   x"D4",   x"82",   x"E3",   x"B5",   x"4F",   x"19", 
  x"F6",   x"A0",   x"5A",   x"0C",   x"6D",   x"3B",   x"C1",   x"97", 
  x"03",   x"55",   x"AF",   x"F9",   x"98",   x"CE",   x"34",   x"62", 
  x"DF",   x"89",   x"73",   x"25",   x"44",   x"12",   x"E8",   x"BE", 
  x"2A",   x"7C",   x"86",   x"D0",   x"B1",   x"E7",   x"1D",   x"4B", 
  x"8B",   x"DD",   x"27",   x"71",   x"10",   x"46",   x"BC",   x"EA", 
  x"7E",   x"28",   x"D2",   x"84",   x"E5",   x"B3",   x"49",   x"1F", 
  x"A2",   x"F4",   x"0E",   x"58",   x"39",   x"6F",   x"95",   x"C3", 
  x"57",   x"01",   x"FB",   x"AD",   x"CC",   x"9A",   x"60",   x"36", 
  x"D9",   x"8F",   x"75",   x"23",   x"42",   x"14",   x"EE",   x"B8", 
  x"2C",   x"7A",   x"80",   x"D6",   x"B7",   x"E1",   x"1B",   x"4D", 
  x"F0",   x"A6",   x"5C",   x"0A",   x"6B",   x"3D",   x"C7",   x"91", 
  x"05",   x"53",   x"A9",   x"FF",   x"9E",   x"C8",   x"32",   x"64", 
  x"2F",   x"79",   x"83",   x"D5",   x"B4",   x"E2",   x"18",   x"4E", 
  x"DA",   x"8C",   x"76",   x"20",   x"41",   x"17",   x"ED",   x"BB", 
  x"06",   x"50",   x"AA",   x"FC",   x"9D",   x"CB",   x"31",   x"67", 
  x"F3",   x"A5",   x"5F",   x"09",   x"68",   x"3E",   x"C4",   x"92", 
  x"7D",   x"2B",   x"D1",   x"87",   x"E6",   x"B0",   x"4A",   x"1C", 
  x"88",   x"DE",   x"24",   x"72",   x"13",   x"45",   x"BF",   x"E9", 
  x"54",   x"02",   x"F8",   x"AE",   x"CF",   x"99",   x"63",   x"35", 
  x"A1",   x"F7",   x"0D",   x"5B",   x"3A",   x"6C",   x"96",   x"C0", 
  x"00",   x"57",   x"AE",   x"F9",   x"9F",   x"C8",   x"31",   x"66", 
  x"FD",   x"AA",   x"53",   x"04",   x"62",   x"35",   x"CC",   x"9B", 
  x"39",   x"6E",   x"97",   x"C0",   x"A6",   x"F1",   x"08",   x"5F", 
  x"C4",   x"93",   x"6A",   x"3D",   x"5B",   x"0C",   x"F5",   x"A2", 
  x"72",   x"25",   x"DC",   x"8B",   x"ED",   x"BA",   x"43",   x"14", 
  x"8F",   x"D8",   x"21",   x"76",   x"10",   x"47",   x"BE",   x"E9", 
  x"4B",   x"1C",   x"E5",   x"B2",   x"D4",   x"83",   x"7A",   x"2D", 
  x"B6",   x"E1",   x"18",   x"4F",   x"29",   x"7E",   x"87",   x"D0", 
  x"E4",   x"B3",   x"4A",   x"1D",   x"7B",   x"2C",   x"D5",   x"82", 
  x"19",   x"4E",   x"B7",   x"E0",   x"86",   x"D1",   x"28",   x"7F", 
  x"DD",   x"8A",   x"73",   x"24",   x"42",   x"15",   x"EC",   x"BB", 
  x"20",   x"77",   x"8E",   x"D9",   x"BF",   x"E8",   x"11",   x"46", 
  x"96",   x"C1",   x"38",   x"6F",   x"09",   x"5E",   x"A7",   x"F0", 
  x"6B",   x"3C",   x"C5",   x"92",   x"F4",   x"A3",   x"5A",   x"0D", 
  x"AF",   x"F8",   x"01",   x"56",   x"30",   x"67",   x"9E",   x"C9", 
  x"52",   x"05",   x"FC",   x"AB",   x"CD",   x"9A",   x"63",   x"34", 
  x"0B",   x"5C",   x"A5",   x"F2",   x"94",   x"C3",   x"3A",   x"6D", 
  x"F6",   x"A1",   x"58",   x"0F",   x"69",   x"3E",   x"C7",   x"90", 
  x"32",   x"65",   x"9C",   x"CB",   x"AD",   x"FA",   x"03",   x"54", 
  x"CF",   x"98",   x"61",   x"36",   x"50",   x"07",   x"FE",   x"A9", 
  x"79",   x"2E",   x"D7",   x"80",   x"E6",   x"B1",   x"48",   x"1F", 
  x"84",   x"D3",   x"2A",   x"7D",   x"1B",   x"4C",   x"B5",   x"E2", 
  x"40",   x"17",   x"EE",   x"B9",   x"DF",   x"88",   x"71",   x"26", 
  x"BD",   x"EA",   x"13",   x"44",   x"22",   x"75",   x"8C",   x"DB", 
  x"EF",   x"B8",   x"41",   x"16",   x"70",   x"27",   x"DE",   x"89", 
  x"12",   x"45",   x"BC",   x"EB",   x"8D",   x"DA",   x"23",   x"74", 
  x"D6",   x"81",   x"78",   x"2F",   x"49",   x"1E",   x"E7",   x"B0", 
  x"2B",   x"7C",   x"85",   x"D2",   x"B4",   x"E3",   x"1A",   x"4D", 
  x"9D",   x"CA",   x"33",   x"64",   x"02",   x"55",   x"AC",   x"FB", 
  x"60",   x"37",   x"CE",   x"99",   x"FF",   x"A8",   x"51",   x"06", 
  x"A4",   x"F3",   x"0A",   x"5D",   x"3B",   x"6C",   x"95",   x"C2", 
  x"59",   x"0E",   x"F7",   x"A0",   x"C6",   x"91",   x"68",   x"3F", 
  x"00",   x"58",   x"B0",   x"E8",   x"A3",   x"FB",   x"13",   x"4B", 
  x"85",   x"DD",   x"35",   x"6D",   x"26",   x"7E",   x"96",   x"CE", 
  x"C9",   x"91",   x"79",   x"21",   x"6A",   x"32",   x"DA",   x"82", 
  x"4C",   x"14",   x"FC",   x"A4",   x"EF",   x"B7",   x"5F",   x"07", 
  x"51",   x"09",   x"E1",   x"B9",   x"F2",   x"AA",   x"42",   x"1A", 
  x"D4",   x"8C",   x"64",   x"3C",   x"77",   x"2F",   x"C7",   x"9F", 
  x"98",   x"C0",   x"28",   x"70",   x"3B",   x"63",   x"8B",   x"D3", 
  x"1D",   x"45",   x"AD",   x"F5",   x"BE",   x"E6",   x"0E",   x"56", 
  x"A2",   x"FA",   x"12",   x"4A",   x"01",   x"59",   x"B1",   x"E9", 
  x"27",   x"7F",   x"97",   x"CF",   x"84",   x"DC",   x"34",   x"6C", 
  x"6B",   x"33",   x"DB",   x"83",   x"C8",   x"90",   x"78",   x"20", 
  x"EE",   x"B6",   x"5E",   x"06",   x"4D",   x"15",   x"FD",   x"A5", 
  x"F3",   x"AB",   x"43",   x"1B",   x"50",   x"08",   x"E0",   x"B8", 
  x"76",   x"2E",   x"C6",   x"9E",   x"D5",   x"8D",   x"65",   x"3D", 
  x"3A",   x"62",   x"8A",   x"D2",   x"99",   x"C1",   x"29",   x"71", 
  x"BF",   x"E7",   x"0F",   x"57",   x"1C",   x"44",   x"AC",   x"F4", 
  x"87",   x"DF",   x"37",   x"6F",   x"24",   x"7C",   x"94",   x"CC", 
  x"02",   x"5A",   x"B2",   x"EA",   x"A1",   x"F9",   x"11",   x"49", 
  x"4E",   x"16",   x"FE",   x"A6",   x"ED",   x"B5",   x"5D",   x"05", 
  x"CB",   x"93",   x"7B",   x"23",   x"68",   x"30",   x"D8",   x"80", 
  x"D6",   x"8E",   x"66",   x"3E",   x"75",   x"2D",   x"C5",   x"9D", 
  x"53",   x"0B",   x"E3",   x"BB",   x"F0",   x"A8",   x"40",   x"18", 
  x"1F",   x"47",   x"AF",   x"F7",   x"BC",   x"E4",   x"0C",   x"54", 
  x"9A",   x"C2",   x"2A",   x"72",   x"39",   x"61",   x"89",   x"D1", 
  x"25",   x"7D",   x"95",   x"CD",   x"86",   x"DE",   x"36",   x"6E", 
  x"A0",   x"F8",   x"10",   x"48",   x"03",   x"5B",   x"B3",   x"EB", 
  x"EC",   x"B4",   x"5C",   x"04",   x"4F",   x"17",   x"FF",   x"A7", 
  x"69",   x"31",   x"D9",   x"81",   x"CA",   x"92",   x"7A",   x"22", 
  x"74",   x"2C",   x"C4",   x"9C",   x"D7",   x"8F",   x"67",   x"3F", 
  x"F1",   x"A9",   x"41",   x"19",   x"52",   x"0A",   x"E2",   x"BA", 
  x"BD",   x"E5",   x"0D",   x"55",   x"1E",   x"46",   x"AE",   x"F6", 
  x"38",   x"60",   x"88",   x"D0",   x"9B",   x"C3",   x"2B",   x"73", 
  x"00",   x"59",   x"B2",   x"EB",   x"A7",   x"FE",   x"15",   x"4C", 
  x"8D",   x"D4",   x"3F",   x"66",   x"2A",   x"73",   x"98",   x"C1", 
  x"D9",   x"80",   x"6B",   x"32",   x"7E",   x"27",   x"CC",   x"95", 
  x"54",   x"0D",   x"E6",   x"BF",   x"F3",   x"AA",   x"41",   x"18", 
  x"71",   x"28",   x"C3",   x"9A",   x"D6",   x"8F",   x"64",   x"3D", 
  x"FC",   x"A5",   x"4E",   x"17",   x"5B",   x"02",   x"E9",   x"B0", 
  x"A8",   x"F1",   x"1A",   x"43",   x"0F",   x"56",   x"BD",   x"E4", 
  x"25",   x"7C",   x"97",   x"CE",   x"82",   x"DB",   x"30",   x"69", 
  x"E2",   x"BB",   x"50",   x"09",   x"45",   x"1C",   x"F7",   x"AE", 
  x"6F",   x"36",   x"DD",   x"84",   x"C8",   x"91",   x"7A",   x"23", 
  x"3B",   x"62",   x"89",   x"D0",   x"9C",   x"C5",   x"2E",   x"77", 
  x"B6",   x"EF",   x"04",   x"5D",   x"11",   x"48",   x"A3",   x"FA", 
  x"93",   x"CA",   x"21",   x"78",   x"34",   x"6D",   x"86",   x"DF", 
  x"1E",   x"47",   x"AC",   x"F5",   x"B9",   x"E0",   x"0B",   x"52", 
  x"4A",   x"13",   x"F8",   x"A1",   x"ED",   x"B4",   x"5F",   x"06", 
  x"C7",   x"9E",   x"75",   x"2C",   x"60",   x"39",   x"D2",   x"8B", 
  x"07",   x"5E",   x"B5",   x"EC",   x"A0",   x"F9",   x"12",   x"4B", 
  x"8A",   x"D3",   x"38",   x"61",   x"2D",   x"74",   x"9F",   x"C6", 
  x"DE",   x"87",   x"6C",   x"35",   x"79",   x"20",   x"CB",   x"92", 
  x"53",   x"0A",   x"E1",   x"B8",   x"F4",   x"AD",   x"46",   x"1F", 
  x"76",   x"2F",   x"C4",   x"9D",   x"D1",   x"88",   x"63",   x"3A", 
  x"FB",   x"A2",   x"49",   x"10",   x"5C",   x"05",   x"EE",   x"B7", 
  x"AF",   x"F6",   x"1D",   x"44",   x"08",   x"51",   x"BA",   x"E3", 
  x"22",   x"7B",   x"90",   x"C9",   x"85",   x"DC",   x"37",   x"6E", 
  x"E5",   x"BC",   x"57",   x"0E",   x"42",   x"1B",   x"F0",   x"A9", 
  x"68",   x"31",   x"DA",   x"83",   x"CF",   x"96",   x"7D",   x"24", 
  x"3C",   x"65",   x"8E",   x"D7",   x"9B",   x"C2",   x"29",   x"70", 
  x"B1",   x"E8",   x"03",   x"5A",   x"16",   x"4F",   x"A4",   x"FD", 
  x"94",   x"CD",   x"26",   x"7F",   x"33",   x"6A",   x"81",   x"D8", 
  x"19",   x"40",   x"AB",   x"F2",   x"BE",   x"E7",   x"0C",   x"55", 
  x"4D",   x"14",   x"FF",   x"A6",   x"EA",   x"B3",   x"58",   x"01", 
  x"C0",   x"99",   x"72",   x"2B",   x"67",   x"3E",   x"D5",   x"8C", 
  x"00",   x"5A",   x"B4",   x"EE",   x"AB",   x"F1",   x"1F",   x"45", 
  x"95",   x"CF",   x"21",   x"7B",   x"3E",   x"64",   x"8A",   x"D0", 
  x"E9",   x"B3",   x"5D",   x"07",   x"42",   x"18",   x"F6",   x"AC", 
  x"7C",   x"26",   x"C8",   x"92",   x"D7",   x"8D",   x"63",   x"39", 
  x"11",   x"4B",   x"A5",   x"FF",   x"BA",   x"E0",   x"0E",   x"54", 
  x"84",   x"DE",   x"30",   x"6A",   x"2F",   x"75",   x"9B",   x"C1", 
  x"F8",   x"A2",   x"4C",   x"16",   x"53",   x"09",   x"E7",   x"BD", 
  x"6D",   x"37",   x"D9",   x"83",   x"C6",   x"9C",   x"72",   x"28", 
  x"22",   x"78",   x"96",   x"CC",   x"89",   x"D3",   x"3D",   x"67", 
  x"B7",   x"ED",   x"03",   x"59",   x"1C",   x"46",   x"A8",   x"F2", 
  x"CB",   x"91",   x"7F",   x"25",   x"60",   x"3A",   x"D4",   x"8E", 
  x"5E",   x"04",   x"EA",   x"B0",   x"F5",   x"AF",   x"41",   x"1B", 
  x"33",   x"69",   x"87",   x"DD",   x"98",   x"C2",   x"2C",   x"76", 
  x"A6",   x"FC",   x"12",   x"48",   x"0D",   x"57",   x"B9",   x"E3", 
  x"DA",   x"80",   x"6E",   x"34",   x"71",   x"2B",   x"C5",   x"9F", 
  x"4F",   x"15",   x"FB",   x"A1",   x"E4",   x"BE",   x"50",   x"0A", 
  x"44",   x"1E",   x"F0",   x"AA",   x"EF",   x"B5",   x"5B",   x"01", 
  x"D1",   x"8B",   x"65",   x"3F",   x"7A",   x"20",   x"CE",   x"94", 
  x"AD",   x"F7",   x"19",   x"43",   x"06",   x"5C",   x"B2",   x"E8", 
  x"38",   x"62",   x"8C",   x"D6",   x"93",   x"C9",   x"27",   x"7D", 
  x"55",   x"0F",   x"E1",   x"BB",   x"FE",   x"A4",   x"4A",   x"10", 
  x"C0",   x"9A",   x"74",   x"2E",   x"6B",   x"31",   x"DF",   x"85", 
  x"BC",   x"E6",   x"08",   x"52",   x"17",   x"4D",   x"A3",   x"F9", 
  x"29",   x"73",   x"9D",   x"C7",   x"82",   x"D8",   x"36",   x"6C", 
  x"66",   x"3C",   x"D2",   x"88",   x"CD",   x"97",   x"79",   x"23", 
  x"F3",   x"A9",   x"47",   x"1D",   x"58",   x"02",   x"EC",   x"B6", 
  x"8F",   x"D5",   x"3B",   x"61",   x"24",   x"7E",   x"90",   x"CA", 
  x"1A",   x"40",   x"AE",   x"F4",   x"B1",   x"EB",   x"05",   x"5F", 
  x"77",   x"2D",   x"C3",   x"99",   x"DC",   x"86",   x"68",   x"32", 
  x"E2",   x"B8",   x"56",   x"0C",   x"49",   x"13",   x"FD",   x"A7", 
  x"9E",   x"C4",   x"2A",   x"70",   x"35",   x"6F",   x"81",   x"DB", 
  x"0B",   x"51",   x"BF",   x"E5",   x"A0",   x"FA",   x"14",   x"4E", 
  x"00",   x"5B",   x"B6",   x"ED",   x"AF",   x"F4",   x"19",   x"42", 
  x"9D",   x"C6",   x"2B",   x"70",   x"32",   x"69",   x"84",   x"DF", 
  x"F9",   x"A2",   x"4F",   x"14",   x"56",   x"0D",   x"E0",   x"BB", 
  x"64",   x"3F",   x"D2",   x"89",   x"CB",   x"90",   x"7D",   x"26", 
  x"31",   x"6A",   x"87",   x"DC",   x"9E",   x"C5",   x"28",   x"73", 
  x"AC",   x"F7",   x"1A",   x"41",   x"03",   x"58",   x"B5",   x"EE", 
  x"C8",   x"93",   x"7E",   x"25",   x"67",   x"3C",   x"D1",   x"8A", 
  x"55",   x"0E",   x"E3",   x"B8",   x"FA",   x"A1",   x"4C",   x"17", 
  x"62",   x"39",   x"D4",   x"8F",   x"CD",   x"96",   x"7B",   x"20", 
  x"FF",   x"A4",   x"49",   x"12",   x"50",   x"0B",   x"E6",   x"BD", 
  x"9B",   x"C0",   x"2D",   x"76",   x"34",   x"6F",   x"82",   x"D9", 
  x"06",   x"5D",   x"B0",   x"EB",   x"A9",   x"F2",   x"1F",   x"44", 
  x"53",   x"08",   x"E5",   x"BE",   x"FC",   x"A7",   x"4A",   x"11", 
  x"CE",   x"95",   x"78",   x"23",   x"61",   x"3A",   x"D7",   x"8C", 
  x"AA",   x"F1",   x"1C",   x"47",   x"05",   x"5E",   x"B3",   x"E8", 
  x"37",   x"6C",   x"81",   x"DA",   x"98",   x"C3",   x"2E",   x"75", 
  x"C4",   x"9F",   x"72",   x"29",   x"6B",   x"30",   x"DD",   x"86", 
  x"59",   x"02",   x"EF",   x"B4",   x"F6",   x"AD",   x"40",   x"1B", 
  x"3D",   x"66",   x"8B",   x"D0",   x"92",   x"C9",   x"24",   x"7F", 
  x"A0",   x"FB",   x"16",   x"4D",   x"0F",   x"54",   x"B9",   x"E2", 
  x"F5",   x"AE",   x"43",   x"18",   x"5A",   x"01",   x"EC",   x"B7", 
  x"68",   x"33",   x"DE",   x"85",   x"C7",   x"9C",   x"71",   x"2A", 
  x"0C",   x"57",   x"BA",   x"E1",   x"A3",   x"F8",   x"15",   x"4E", 
  x"91",   x"CA",   x"27",   x"7C",   x"3E",   x"65",   x"88",   x"D3", 
  x"A6",   x"FD",   x"10",   x"4B",   x"09",   x"52",   x"BF",   x"E4", 
  x"3B",   x"60",   x"8D",   x"D6",   x"94",   x"CF",   x"22",   x"79", 
  x"5F",   x"04",   x"E9",   x"B2",   x"F0",   x"AB",   x"46",   x"1D", 
  x"C2",   x"99",   x"74",   x"2F",   x"6D",   x"36",   x"DB",   x"80", 
  x"97",   x"CC",   x"21",   x"7A",   x"38",   x"63",   x"8E",   x"D5", 
  x"0A",   x"51",   x"BC",   x"E7",   x"A5",   x"FE",   x"13",   x"48", 
  x"6E",   x"35",   x"D8",   x"83",   x"C1",   x"9A",   x"77",   x"2C", 
  x"F3",   x"A8",   x"45",   x"1E",   x"5C",   x"07",   x"EA",   x"B1", 
  x"00",   x"5C",   x"B8",   x"E4",   x"B3",   x"EF",   x"0B",   x"57", 
  x"A5",   x"F9",   x"1D",   x"41",   x"16",   x"4A",   x"AE",   x"F2", 
  x"89",   x"D5",   x"31",   x"6D",   x"3A",   x"66",   x"82",   x"DE", 
  x"2C",   x"70",   x"94",   x"C8",   x"9F",   x"C3",   x"27",   x"7B", 
  x"D1",   x"8D",   x"69",   x"35",   x"62",   x"3E",   x"DA",   x"86", 
  x"74",   x"28",   x"CC",   x"90",   x"C7",   x"9B",   x"7F",   x"23", 
  x"58",   x"04",   x"E0",   x"BC",   x"EB",   x"B7",   x"53",   x"0F", 
  x"FD",   x"A1",   x"45",   x"19",   x"4E",   x"12",   x"F6",   x"AA", 
  x"61",   x"3D",   x"D9",   x"85",   x"D2",   x"8E",   x"6A",   x"36", 
  x"C4",   x"98",   x"7C",   x"20",   x"77",   x"2B",   x"CF",   x"93", 
  x"E8",   x"B4",   x"50",   x"0C",   x"5B",   x"07",   x"E3",   x"BF", 
  x"4D",   x"11",   x"F5",   x"A9",   x"FE",   x"A2",   x"46",   x"1A", 
  x"B0",   x"EC",   x"08",   x"54",   x"03",   x"5F",   x"BB",   x"E7", 
  x"15",   x"49",   x"AD",   x"F1",   x"A6",   x"FA",   x"1E",   x"42", 
  x"39",   x"65",   x"81",   x"DD",   x"8A",   x"D6",   x"32",   x"6E", 
  x"9C",   x"C0",   x"24",   x"78",   x"2F",   x"73",   x"97",   x"CB", 
  x"C2",   x"9E",   x"7A",   x"26",   x"71",   x"2D",   x"C9",   x"95", 
  x"67",   x"3B",   x"DF",   x"83",   x"D4",   x"88",   x"6C",   x"30", 
  x"4B",   x"17",   x"F3",   x"AF",   x"F8",   x"A4",   x"40",   x"1C", 
  x"EE",   x"B2",   x"56",   x"0A",   x"5D",   x"01",   x"E5",   x"B9", 
  x"13",   x"4F",   x"AB",   x"F7",   x"A0",   x"FC",   x"18",   x"44", 
  x"B6",   x"EA",   x"0E",   x"52",   x"05",   x"59",   x"BD",   x"E1", 
  x"9A",   x"C6",   x"22",   x"7E",   x"29",   x"75",   x"91",   x"CD", 
  x"3F",   x"63",   x"87",   x"DB",   x"8C",   x"D0",   x"34",   x"68", 
  x"A3",   x"FF",   x"1B",   x"47",   x"10",   x"4C",   x"A8",   x"F4", 
  x"06",   x"5A",   x"BE",   x"E2",   x"B5",   x"E9",   x"0D",   x"51", 
  x"2A",   x"76",   x"92",   x"CE",   x"99",   x"C5",   x"21",   x"7D", 
  x"8F",   x"D3",   x"37",   x"6B",   x"3C",   x"60",   x"84",   x"D8", 
  x"72",   x"2E",   x"CA",   x"96",   x"C1",   x"9D",   x"79",   x"25", 
  x"D7",   x"8B",   x"6F",   x"33",   x"64",   x"38",   x"DC",   x"80", 
  x"FB",   x"A7",   x"43",   x"1F",   x"48",   x"14",   x"F0",   x"AC", 
  x"5E",   x"02",   x"E6",   x"BA",   x"ED",   x"B1",   x"55",   x"09", 
  x"00",   x"5D",   x"BA",   x"E7",   x"B7",   x"EA",   x"0D",   x"50", 
  x"AD",   x"F0",   x"17",   x"4A",   x"1A",   x"47",   x"A0",   x"FD", 
  x"99",   x"C4",   x"23",   x"7E",   x"2E",   x"73",   x"94",   x"C9", 
  x"34",   x"69",   x"8E",   x"D3",   x"83",   x"DE",   x"39",   x"64", 
  x"F1",   x"AC",   x"4B",   x"16",   x"46",   x"1B",   x"FC",   x"A1", 
  x"5C",   x"01",   x"E6",   x"BB",   x"EB",   x"B6",   x"51",   x"0C", 
  x"68",   x"35",   x"D2",   x"8F",   x"DF",   x"82",   x"65",   x"38", 
  x"C5",   x"98",   x"7F",   x"22",   x"72",   x"2F",   x"C8",   x"95", 
  x"21",   x"7C",   x"9B",   x"C6",   x"96",   x"CB",   x"2C",   x"71", 
  x"8C",   x"D1",   x"36",   x"6B",   x"3B",   x"66",   x"81",   x"DC", 
  x"B8",   x"E5",   x"02",   x"5F",   x"0F",   x"52",   x"B5",   x"E8", 
  x"15",   x"48",   x"AF",   x"F2",   x"A2",   x"FF",   x"18",   x"45", 
  x"D0",   x"8D",   x"6A",   x"37",   x"67",   x"3A",   x"DD",   x"80", 
  x"7D",   x"20",   x"C7",   x"9A",   x"CA",   x"97",   x"70",   x"2D", 
  x"49",   x"14",   x"F3",   x"AE",   x"FE",   x"A3",   x"44",   x"19", 
  x"E4",   x"B9",   x"5E",   x"03",   x"53",   x"0E",   x"E9",   x"B4", 
  x"42",   x"1F",   x"F8",   x"A5",   x"F5",   x"A8",   x"4F",   x"12", 
  x"EF",   x"B2",   x"55",   x"08",   x"58",   x"05",   x"E2",   x"BF", 
  x"DB",   x"86",   x"61",   x"3C",   x"6C",   x"31",   x"D6",   x"8B", 
  x"76",   x"2B",   x"CC",   x"91",   x"C1",   x"9C",   x"7B",   x"26", 
  x"B3",   x"EE",   x"09",   x"54",   x"04",   x"59",   x"BE",   x"E3", 
  x"1E",   x"43",   x"A4",   x"F9",   x"A9",   x"F4",   x"13",   x"4E", 
  x"2A",   x"77",   x"90",   x"CD",   x"9D",   x"C0",   x"27",   x"7A", 
  x"87",   x"DA",   x"3D",   x"60",   x"30",   x"6D",   x"8A",   x"D7", 
  x"63",   x"3E",   x"D9",   x"84",   x"D4",   x"89",   x"6E",   x"33", 
  x"CE",   x"93",   x"74",   x"29",   x"79",   x"24",   x"C3",   x"9E", 
  x"FA",   x"A7",   x"40",   x"1D",   x"4D",   x"10",   x"F7",   x"AA", 
  x"57",   x"0A",   x"ED",   x"B0",   x"E0",   x"BD",   x"5A",   x"07", 
  x"92",   x"CF",   x"28",   x"75",   x"25",   x"78",   x"9F",   x"C2", 
  x"3F",   x"62",   x"85",   x"D8",   x"88",   x"D5",   x"32",   x"6F", 
  x"0B",   x"56",   x"B1",   x"EC",   x"BC",   x"E1",   x"06",   x"5B", 
  x"A6",   x"FB",   x"1C",   x"41",   x"11",   x"4C",   x"AB",   x"F6", 
  x"00",   x"5E",   x"BC",   x"E2",   x"BB",   x"E5",   x"07",   x"59", 
  x"B5",   x"EB",   x"09",   x"57",   x"0E",   x"50",   x"B2",   x"EC", 
  x"A9",   x"F7",   x"15",   x"4B",   x"12",   x"4C",   x"AE",   x"F0", 
  x"1C",   x"42",   x"A0",   x"FE",   x"A7",   x"F9",   x"1B",   x"45", 
  x"91",   x"CF",   x"2D",   x"73",   x"2A",   x"74",   x"96",   x"C8", 
  x"24",   x"7A",   x"98",   x"C6",   x"9F",   x"C1",   x"23",   x"7D", 
  x"38",   x"66",   x"84",   x"DA",   x"83",   x"DD",   x"3F",   x"61", 
  x"8D",   x"D3",   x"31",   x"6F",   x"36",   x"68",   x"8A",   x"D4", 
  x"E1",   x"BF",   x"5D",   x"03",   x"5A",   x"04",   x"E6",   x"B8", 
  x"54",   x"0A",   x"E8",   x"B6",   x"EF",   x"B1",   x"53",   x"0D", 
  x"48",   x"16",   x"F4",   x"AA",   x"F3",   x"AD",   x"4F",   x"11", 
  x"FD",   x"A3",   x"41",   x"1F",   x"46",   x"18",   x"FA",   x"A4", 
  x"70",   x"2E",   x"CC",   x"92",   x"CB",   x"95",   x"77",   x"29", 
  x"C5",   x"9B",   x"79",   x"27",   x"7E",   x"20",   x"C2",   x"9C", 
  x"D9",   x"87",   x"65",   x"3B",   x"62",   x"3C",   x"DE",   x"80", 
  x"6C",   x"32",   x"D0",   x"8E",   x"D7",   x"89",   x"6B",   x"35", 
  x"01",   x"5F",   x"BD",   x"E3",   x"BA",   x"E4",   x"06",   x"58", 
  x"B4",   x"EA",   x"08",   x"56",   x"0F",   x"51",   x"B3",   x"ED", 
  x"A8",   x"F6",   x"14",   x"4A",   x"13",   x"4D",   x"AF",   x"F1", 
  x"1D",   x"43",   x"A1",   x"FF",   x"A6",   x"F8",   x"1A",   x"44", 
  x"90",   x"CE",   x"2C",   x"72",   x"2B",   x"75",   x"97",   x"C9", 
  x"25",   x"7B",   x"99",   x"C7",   x"9E",   x"C0",   x"22",   x"7C", 
  x"39",   x"67",   x"85",   x"DB",   x"82",   x"DC",   x"3E",   x"60", 
  x"8C",   x"D2",   x"30",   x"6E",   x"37",   x"69",   x"8B",   x"D5", 
  x"E0",   x"BE",   x"5C",   x"02",   x"5B",   x"05",   x"E7",   x"B9", 
  x"55",   x"0B",   x"E9",   x"B7",   x"EE",   x"B0",   x"52",   x"0C", 
  x"49",   x"17",   x"F5",   x"AB",   x"F2",   x"AC",   x"4E",   x"10", 
  x"FC",   x"A2",   x"40",   x"1E",   x"47",   x"19",   x"FB",   x"A5", 
  x"71",   x"2F",   x"CD",   x"93",   x"CA",   x"94",   x"76",   x"28", 
  x"C4",   x"9A",   x"78",   x"26",   x"7F",   x"21",   x"C3",   x"9D", 
  x"D8",   x"86",   x"64",   x"3A",   x"63",   x"3D",   x"DF",   x"81", 
  x"6D",   x"33",   x"D1",   x"8F",   x"D6",   x"88",   x"6A",   x"34", 
  x"00",   x"5F",   x"BE",   x"E1",   x"BF",   x"E0",   x"01",   x"5E", 
  x"BD",   x"E2",   x"03",   x"5C",   x"02",   x"5D",   x"BC",   x"E3", 
  x"B9",   x"E6",   x"07",   x"58",   x"06",   x"59",   x"B8",   x"E7", 
  x"04",   x"5B",   x"BA",   x"E5",   x"BB",   x"E4",   x"05",   x"5A", 
  x"B1",   x"EE",   x"0F",   x"50",   x"0E",   x"51",   x"B0",   x"EF", 
  x"0C",   x"53",   x"B2",   x"ED",   x"B3",   x"EC",   x"0D",   x"52", 
  x"08",   x"57",   x"B6",   x"E9",   x"B7",   x"E8",   x"09",   x"56", 
  x"B5",   x"EA",   x"0B",   x"54",   x"0A",   x"55",   x"B4",   x"EB", 
  x"A1",   x"FE",   x"1F",   x"40",   x"1E",   x"41",   x"A0",   x"FF", 
  x"1C",   x"43",   x"A2",   x"FD",   x"A3",   x"FC",   x"1D",   x"42", 
  x"18",   x"47",   x"A6",   x"F9",   x"A7",   x"F8",   x"19",   x"46", 
  x"A5",   x"FA",   x"1B",   x"44",   x"1A",   x"45",   x"A4",   x"FB", 
  x"10",   x"4F",   x"AE",   x"F1",   x"AF",   x"F0",   x"11",   x"4E", 
  x"AD",   x"F2",   x"13",   x"4C",   x"12",   x"4D",   x"AC",   x"F3", 
  x"A9",   x"F6",   x"17",   x"48",   x"16",   x"49",   x"A8",   x"F7", 
  x"14",   x"4B",   x"AA",   x"F5",   x"AB",   x"F4",   x"15",   x"4A", 
  x"81",   x"DE",   x"3F",   x"60",   x"3E",   x"61",   x"80",   x"DF", 
  x"3C",   x"63",   x"82",   x"DD",   x"83",   x"DC",   x"3D",   x"62", 
  x"38",   x"67",   x"86",   x"D9",   x"87",   x"D8",   x"39",   x"66", 
  x"85",   x"DA",   x"3B",   x"64",   x"3A",   x"65",   x"84",   x"DB", 
  x"30",   x"6F",   x"8E",   x"D1",   x"8F",   x"D0",   x"31",   x"6E", 
  x"8D",   x"D2",   x"33",   x"6C",   x"32",   x"6D",   x"8C",   x"D3", 
  x"89",   x"D6",   x"37",   x"68",   x"36",   x"69",   x"88",   x"D7", 
  x"34",   x"6B",   x"8A",   x"D5",   x"8B",   x"D4",   x"35",   x"6A", 
  x"20",   x"7F",   x"9E",   x"C1",   x"9F",   x"C0",   x"21",   x"7E", 
  x"9D",   x"C2",   x"23",   x"7C",   x"22",   x"7D",   x"9C",   x"C3", 
  x"99",   x"C6",   x"27",   x"78",   x"26",   x"79",   x"98",   x"C7", 
  x"24",   x"7B",   x"9A",   x"C5",   x"9B",   x"C4",   x"25",   x"7A", 
  x"91",   x"CE",   x"2F",   x"70",   x"2E",   x"71",   x"90",   x"CF", 
  x"2C",   x"73",   x"92",   x"CD",   x"93",   x"CC",   x"2D",   x"72", 
  x"28",   x"77",   x"96",   x"C9",   x"97",   x"C8",   x"29",   x"76", 
  x"95",   x"CA",   x"2B",   x"74",   x"2A",   x"75",   x"94",   x"CB", 
  x"00",   x"60",   x"C0",   x"A0",   x"43",   x"23",   x"83",   x"E3", 
  x"86",   x"E6",   x"46",   x"26",   x"C5",   x"A5",   x"05",   x"65", 
  x"CF",   x"AF",   x"0F",   x"6F",   x"8C",   x"EC",   x"4C",   x"2C", 
  x"49",   x"29",   x"89",   x"E9",   x"0A",   x"6A",   x"CA",   x"AA", 
  x"5D",   x"3D",   x"9D",   x"FD",   x"1E",   x"7E",   x"DE",   x"BE", 
  x"DB",   x"BB",   x"1B",   x"7B",   x"98",   x"F8",   x"58",   x"38", 
  x"92",   x"F2",   x"52",   x"32",   x"D1",   x"B1",   x"11",   x"71", 
  x"14",   x"74",   x"D4",   x"B4",   x"57",   x"37",   x"97",   x"F7", 
  x"BA",   x"DA",   x"7A",   x"1A",   x"F9",   x"99",   x"39",   x"59", 
  x"3C",   x"5C",   x"FC",   x"9C",   x"7F",   x"1F",   x"BF",   x"DF", 
  x"75",   x"15",   x"B5",   x"D5",   x"36",   x"56",   x"F6",   x"96", 
  x"F3",   x"93",   x"33",   x"53",   x"B0",   x"D0",   x"70",   x"10", 
  x"E7",   x"87",   x"27",   x"47",   x"A4",   x"C4",   x"64",   x"04", 
  x"61",   x"01",   x"A1",   x"C1",   x"22",   x"42",   x"E2",   x"82", 
  x"28",   x"48",   x"E8",   x"88",   x"6B",   x"0B",   x"AB",   x"CB", 
  x"AE",   x"CE",   x"6E",   x"0E",   x"ED",   x"8D",   x"2D",   x"4D", 
  x"B7",   x"D7",   x"77",   x"17",   x"F4",   x"94",   x"34",   x"54", 
  x"31",   x"51",   x"F1",   x"91",   x"72",   x"12",   x"B2",   x"D2", 
  x"78",   x"18",   x"B8",   x"D8",   x"3B",   x"5B",   x"FB",   x"9B", 
  x"FE",   x"9E",   x"3E",   x"5E",   x"BD",   x"DD",   x"7D",   x"1D", 
  x"EA",   x"8A",   x"2A",   x"4A",   x"A9",   x"C9",   x"69",   x"09", 
  x"6C",   x"0C",   x"AC",   x"CC",   x"2F",   x"4F",   x"EF",   x"8F", 
  x"25",   x"45",   x"E5",   x"85",   x"66",   x"06",   x"A6",   x"C6", 
  x"A3",   x"C3",   x"63",   x"03",   x"E0",   x"80",   x"20",   x"40", 
  x"0D",   x"6D",   x"CD",   x"AD",   x"4E",   x"2E",   x"8E",   x"EE", 
  x"8B",   x"EB",   x"4B",   x"2B",   x"C8",   x"A8",   x"08",   x"68", 
  x"C2",   x"A2",   x"02",   x"62",   x"81",   x"E1",   x"41",   x"21", 
  x"44",   x"24",   x"84",   x"E4",   x"07",   x"67",   x"C7",   x"A7", 
  x"50",   x"30",   x"90",   x"F0",   x"13",   x"73",   x"D3",   x"B3", 
  x"D6",   x"B6",   x"16",   x"76",   x"95",   x"F5",   x"55",   x"35", 
  x"9F",   x"FF",   x"5F",   x"3F",   x"DC",   x"BC",   x"1C",   x"7C", 
  x"19",   x"79",   x"D9",   x"B9",   x"5A",   x"3A",   x"9A",   x"FA", 
  x"00",   x"61",   x"C2",   x"A3",   x"47",   x"26",   x"85",   x"E4", 
  x"8E",   x"EF",   x"4C",   x"2D",   x"C9",   x"A8",   x"0B",   x"6A", 
  x"DF",   x"BE",   x"1D",   x"7C",   x"98",   x"F9",   x"5A",   x"3B", 
  x"51",   x"30",   x"93",   x"F2",   x"16",   x"77",   x"D4",   x"B5", 
  x"7D",   x"1C",   x"BF",   x"DE",   x"3A",   x"5B",   x"F8",   x"99", 
  x"F3",   x"92",   x"31",   x"50",   x"B4",   x"D5",   x"76",   x"17", 
  x"A2",   x"C3",   x"60",   x"01",   x"E5",   x"84",   x"27",   x"46", 
  x"2C",   x"4D",   x"EE",   x"8F",   x"6B",   x"0A",   x"A9",   x"C8", 
  x"FA",   x"9B",   x"38",   x"59",   x"BD",   x"DC",   x"7F",   x"1E", 
  x"74",   x"15",   x"B6",   x"D7",   x"33",   x"52",   x"F1",   x"90", 
  x"25",   x"44",   x"E7",   x"86",   x"62",   x"03",   x"A0",   x"C1", 
  x"AB",   x"CA",   x"69",   x"08",   x"EC",   x"8D",   x"2E",   x"4F", 
  x"87",   x"E6",   x"45",   x"24",   x"C0",   x"A1",   x"02",   x"63", 
  x"09",   x"68",   x"CB",   x"AA",   x"4E",   x"2F",   x"8C",   x"ED", 
  x"58",   x"39",   x"9A",   x"FB",   x"1F",   x"7E",   x"DD",   x"BC", 
  x"D6",   x"B7",   x"14",   x"75",   x"91",   x"F0",   x"53",   x"32", 
  x"37",   x"56",   x"F5",   x"94",   x"70",   x"11",   x"B2",   x"D3", 
  x"B9",   x"D8",   x"7B",   x"1A",   x"FE",   x"9F",   x"3C",   x"5D", 
  x"E8",   x"89",   x"2A",   x"4B",   x"AF",   x"CE",   x"6D",   x"0C", 
  x"66",   x"07",   x"A4",   x"C5",   x"21",   x"40",   x"E3",   x"82", 
  x"4A",   x"2B",   x"88",   x"E9",   x"0D",   x"6C",   x"CF",   x"AE", 
  x"C4",   x"A5",   x"06",   x"67",   x"83",   x"E2",   x"41",   x"20", 
  x"95",   x"F4",   x"57",   x"36",   x"D2",   x"B3",   x"10",   x"71", 
  x"1B",   x"7A",   x"D9",   x"B8",   x"5C",   x"3D",   x"9E",   x"FF", 
  x"CD",   x"AC",   x"0F",   x"6E",   x"8A",   x"EB",   x"48",   x"29", 
  x"43",   x"22",   x"81",   x"E0",   x"04",   x"65",   x"C6",   x"A7", 
  x"12",   x"73",   x"D0",   x"B1",   x"55",   x"34",   x"97",   x"F6", 
  x"9C",   x"FD",   x"5E",   x"3F",   x"DB",   x"BA",   x"19",   x"78", 
  x"B0",   x"D1",   x"72",   x"13",   x"F7",   x"96",   x"35",   x"54", 
  x"3E",   x"5F",   x"FC",   x"9D",   x"79",   x"18",   x"BB",   x"DA", 
  x"6F",   x"0E",   x"AD",   x"CC",   x"28",   x"49",   x"EA",   x"8B", 
  x"E1",   x"80",   x"23",   x"42",   x"A6",   x"C7",   x"64",   x"05", 
  x"00",   x"62",   x"C4",   x"A6",   x"4B",   x"29",   x"8F",   x"ED", 
  x"96",   x"F4",   x"52",   x"30",   x"DD",   x"BF",   x"19",   x"7B", 
  x"EF",   x"8D",   x"2B",   x"49",   x"A4",   x"C6",   x"60",   x"02", 
  x"79",   x"1B",   x"BD",   x"DF",   x"32",   x"50",   x"F6",   x"94", 
  x"1D",   x"7F",   x"D9",   x"BB",   x"56",   x"34",   x"92",   x"F0", 
  x"8B",   x"E9",   x"4F",   x"2D",   x"C0",   x"A2",   x"04",   x"66", 
  x"F2",   x"90",   x"36",   x"54",   x"B9",   x"DB",   x"7D",   x"1F", 
  x"64",   x"06",   x"A0",   x"C2",   x"2F",   x"4D",   x"EB",   x"89", 
  x"3A",   x"58",   x"FE",   x"9C",   x"71",   x"13",   x"B5",   x"D7", 
  x"AC",   x"CE",   x"68",   x"0A",   x"E7",   x"85",   x"23",   x"41", 
  x"D5",   x"B7",   x"11",   x"73",   x"9E",   x"FC",   x"5A",   x"38", 
  x"43",   x"21",   x"87",   x"E5",   x"08",   x"6A",   x"CC",   x"AE", 
  x"27",   x"45",   x"E3",   x"81",   x"6C",   x"0E",   x"A8",   x"CA", 
  x"B1",   x"D3",   x"75",   x"17",   x"FA",   x"98",   x"3E",   x"5C", 
  x"C8",   x"AA",   x"0C",   x"6E",   x"83",   x"E1",   x"47",   x"25", 
  x"5E",   x"3C",   x"9A",   x"F8",   x"15",   x"77",   x"D1",   x"B3", 
  x"74",   x"16",   x"B0",   x"D2",   x"3F",   x"5D",   x"FB",   x"99", 
  x"E2",   x"80",   x"26",   x"44",   x"A9",   x"CB",   x"6D",   x"0F", 
  x"9B",   x"F9",   x"5F",   x"3D",   x"D0",   x"B2",   x"14",   x"76", 
  x"0D",   x"6F",   x"C9",   x"AB",   x"46",   x"24",   x"82",   x"E0", 
  x"69",   x"0B",   x"AD",   x"CF",   x"22",   x"40",   x"E6",   x"84", 
  x"FF",   x"9D",   x"3B",   x"59",   x"B4",   x"D6",   x"70",   x"12", 
  x"86",   x"E4",   x"42",   x"20",   x"CD",   x"AF",   x"09",   x"6B", 
  x"10",   x"72",   x"D4",   x"B6",   x"5B",   x"39",   x"9F",   x"FD", 
  x"4E",   x"2C",   x"8A",   x"E8",   x"05",   x"67",   x"C1",   x"A3", 
  x"D8",   x"BA",   x"1C",   x"7E",   x"93",   x"F1",   x"57",   x"35", 
  x"A1",   x"C3",   x"65",   x"07",   x"EA",   x"88",   x"2E",   x"4C", 
  x"37",   x"55",   x"F3",   x"91",   x"7C",   x"1E",   x"B8",   x"DA", 
  x"53",   x"31",   x"97",   x"F5",   x"18",   x"7A",   x"DC",   x"BE", 
  x"C5",   x"A7",   x"01",   x"63",   x"8E",   x"EC",   x"4A",   x"28", 
  x"BC",   x"DE",   x"78",   x"1A",   x"F7",   x"95",   x"33",   x"51", 
  x"2A",   x"48",   x"EE",   x"8C",   x"61",   x"03",   x"A5",   x"C7", 
  x"00",   x"63",   x"C6",   x"A5",   x"4F",   x"2C",   x"89",   x"EA", 
  x"9E",   x"FD",   x"58",   x"3B",   x"D1",   x"B2",   x"17",   x"74", 
  x"FF",   x"9C",   x"39",   x"5A",   x"B0",   x"D3",   x"76",   x"15", 
  x"61",   x"02",   x"A7",   x"C4",   x"2E",   x"4D",   x"E8",   x"8B", 
  x"3D",   x"5E",   x"FB",   x"98",   x"72",   x"11",   x"B4",   x"D7", 
  x"A3",   x"C0",   x"65",   x"06",   x"EC",   x"8F",   x"2A",   x"49", 
  x"C2",   x"A1",   x"04",   x"67",   x"8D",   x"EE",   x"4B",   x"28", 
  x"5C",   x"3F",   x"9A",   x"F9",   x"13",   x"70",   x"D5",   x"B6", 
  x"7A",   x"19",   x"BC",   x"DF",   x"35",   x"56",   x"F3",   x"90", 
  x"E4",   x"87",   x"22",   x"41",   x"AB",   x"C8",   x"6D",   x"0E", 
  x"85",   x"E6",   x"43",   x"20",   x"CA",   x"A9",   x"0C",   x"6F", 
  x"1B",   x"78",   x"DD",   x"BE",   x"54",   x"37",   x"92",   x"F1", 
  x"47",   x"24",   x"81",   x"E2",   x"08",   x"6B",   x"CE",   x"AD", 
  x"D9",   x"BA",   x"1F",   x"7C",   x"96",   x"F5",   x"50",   x"33", 
  x"B8",   x"DB",   x"7E",   x"1D",   x"F7",   x"94",   x"31",   x"52", 
  x"26",   x"45",   x"E0",   x"83",   x"69",   x"0A",   x"AF",   x"CC", 
  x"F4",   x"97",   x"32",   x"51",   x"BB",   x"D8",   x"7D",   x"1E", 
  x"6A",   x"09",   x"AC",   x"CF",   x"25",   x"46",   x"E3",   x"80", 
  x"0B",   x"68",   x"CD",   x"AE",   x"44",   x"27",   x"82",   x"E1", 
  x"95",   x"F6",   x"53",   x"30",   x"DA",   x"B9",   x"1C",   x"7F", 
  x"C9",   x"AA",   x"0F",   x"6C",   x"86",   x"E5",   x"40",   x"23", 
  x"57",   x"34",   x"91",   x"F2",   x"18",   x"7B",   x"DE",   x"BD", 
  x"36",   x"55",   x"F0",   x"93",   x"79",   x"1A",   x"BF",   x"DC", 
  x"A8",   x"CB",   x"6E",   x"0D",   x"E7",   x"84",   x"21",   x"42", 
  x"8E",   x"ED",   x"48",   x"2B",   x"C1",   x"A2",   x"07",   x"64", 
  x"10",   x"73",   x"D6",   x"B5",   x"5F",   x"3C",   x"99",   x"FA", 
  x"71",   x"12",   x"B7",   x"D4",   x"3E",   x"5D",   x"F8",   x"9B", 
  x"EF",   x"8C",   x"29",   x"4A",   x"A0",   x"C3",   x"66",   x"05", 
  x"B3",   x"D0",   x"75",   x"16",   x"FC",   x"9F",   x"3A",   x"59", 
  x"2D",   x"4E",   x"EB",   x"88",   x"62",   x"01",   x"A4",   x"C7", 
  x"4C",   x"2F",   x"8A",   x"E9",   x"03",   x"60",   x"C5",   x"A6", 
  x"D2",   x"B1",   x"14",   x"77",   x"9D",   x"FE",   x"5B",   x"38", 
  x"00",   x"64",   x"C8",   x"AC",   x"53",   x"37",   x"9B",   x"FF", 
  x"A6",   x"C2",   x"6E",   x"0A",   x"F5",   x"91",   x"3D",   x"59", 
  x"8F",   x"EB",   x"47",   x"23",   x"DC",   x"B8",   x"14",   x"70", 
  x"29",   x"4D",   x"E1",   x"85",   x"7A",   x"1E",   x"B2",   x"D6", 
  x"DD",   x"B9",   x"15",   x"71",   x"8E",   x"EA",   x"46",   x"22", 
  x"7B",   x"1F",   x"B3",   x"D7",   x"28",   x"4C",   x"E0",   x"84", 
  x"52",   x"36",   x"9A",   x"FE",   x"01",   x"65",   x"C9",   x"AD", 
  x"F4",   x"90",   x"3C",   x"58",   x"A7",   x"C3",   x"6F",   x"0B", 
  x"79",   x"1D",   x"B1",   x"D5",   x"2A",   x"4E",   x"E2",   x"86", 
  x"DF",   x"BB",   x"17",   x"73",   x"8C",   x"E8",   x"44",   x"20", 
  x"F6",   x"92",   x"3E",   x"5A",   x"A5",   x"C1",   x"6D",   x"09", 
  x"50",   x"34",   x"98",   x"FC",   x"03",   x"67",   x"CB",   x"AF", 
  x"A4",   x"C0",   x"6C",   x"08",   x"F7",   x"93",   x"3F",   x"5B", 
  x"02",   x"66",   x"CA",   x"AE",   x"51",   x"35",   x"99",   x"FD", 
  x"2B",   x"4F",   x"E3",   x"87",   x"78",   x"1C",   x"B0",   x"D4", 
  x"8D",   x"E9",   x"45",   x"21",   x"DE",   x"BA",   x"16",   x"72", 
  x"F2",   x"96",   x"3A",   x"5E",   x"A1",   x"C5",   x"69",   x"0D", 
  x"54",   x"30",   x"9C",   x"F8",   x"07",   x"63",   x"CF",   x"AB", 
  x"7D",   x"19",   x"B5",   x"D1",   x"2E",   x"4A",   x"E6",   x"82", 
  x"DB",   x"BF",   x"13",   x"77",   x"88",   x"EC",   x"40",   x"24", 
  x"2F",   x"4B",   x"E7",   x"83",   x"7C",   x"18",   x"B4",   x"D0", 
  x"89",   x"ED",   x"41",   x"25",   x"DA",   x"BE",   x"12",   x"76", 
  x"A0",   x"C4",   x"68",   x"0C",   x"F3",   x"97",   x"3B",   x"5F", 
  x"06",   x"62",   x"CE",   x"AA",   x"55",   x"31",   x"9D",   x"F9", 
  x"8B",   x"EF",   x"43",   x"27",   x"D8",   x"BC",   x"10",   x"74", 
  x"2D",   x"49",   x"E5",   x"81",   x"7E",   x"1A",   x"B6",   x"D2", 
  x"04",   x"60",   x"CC",   x"A8",   x"57",   x"33",   x"9F",   x"FB", 
  x"A2",   x"C6",   x"6A",   x"0E",   x"F1",   x"95",   x"39",   x"5D", 
  x"56",   x"32",   x"9E",   x"FA",   x"05",   x"61",   x"CD",   x"A9", 
  x"F0",   x"94",   x"38",   x"5C",   x"A3",   x"C7",   x"6B",   x"0F", 
  x"D9",   x"BD",   x"11",   x"75",   x"8A",   x"EE",   x"42",   x"26", 
  x"7F",   x"1B",   x"B7",   x"D3",   x"2C",   x"48",   x"E4",   x"80", 
  x"00",   x"65",   x"CA",   x"AF",   x"57",   x"32",   x"9D",   x"F8", 
  x"AE",   x"CB",   x"64",   x"01",   x"F9",   x"9C",   x"33",   x"56", 
  x"9F",   x"FA",   x"55",   x"30",   x"C8",   x"AD",   x"02",   x"67", 
  x"31",   x"54",   x"FB",   x"9E",   x"66",   x"03",   x"AC",   x"C9", 
  x"FD",   x"98",   x"37",   x"52",   x"AA",   x"CF",   x"60",   x"05", 
  x"53",   x"36",   x"99",   x"FC",   x"04",   x"61",   x"CE",   x"AB", 
  x"62",   x"07",   x"A8",   x"CD",   x"35",   x"50",   x"FF",   x"9A", 
  x"CC",   x"A9",   x"06",   x"63",   x"9B",   x"FE",   x"51",   x"34", 
  x"39",   x"5C",   x"F3",   x"96",   x"6E",   x"0B",   x"A4",   x"C1", 
  x"97",   x"F2",   x"5D",   x"38",   x"C0",   x"A5",   x"0A",   x"6F", 
  x"A6",   x"C3",   x"6C",   x"09",   x"F1",   x"94",   x"3B",   x"5E", 
  x"08",   x"6D",   x"C2",   x"A7",   x"5F",   x"3A",   x"95",   x"F0", 
  x"C4",   x"A1",   x"0E",   x"6B",   x"93",   x"F6",   x"59",   x"3C", 
  x"6A",   x"0F",   x"A0",   x"C5",   x"3D",   x"58",   x"F7",   x"92", 
  x"5B",   x"3E",   x"91",   x"F4",   x"0C",   x"69",   x"C6",   x"A3", 
  x"F5",   x"90",   x"3F",   x"5A",   x"A2",   x"C7",   x"68",   x"0D", 
  x"72",   x"17",   x"B8",   x"DD",   x"25",   x"40",   x"EF",   x"8A", 
  x"DC",   x"B9",   x"16",   x"73",   x"8B",   x"EE",   x"41",   x"24", 
  x"ED",   x"88",   x"27",   x"42",   x"BA",   x"DF",   x"70",   x"15", 
  x"43",   x"26",   x"89",   x"EC",   x"14",   x"71",   x"DE",   x"BB", 
  x"8F",   x"EA",   x"45",   x"20",   x"D8",   x"BD",   x"12",   x"77", 
  x"21",   x"44",   x"EB",   x"8E",   x"76",   x"13",   x"BC",   x"D9", 
  x"10",   x"75",   x"DA",   x"BF",   x"47",   x"22",   x"8D",   x"E8", 
  x"BE",   x"DB",   x"74",   x"11",   x"E9",   x"8C",   x"23",   x"46", 
  x"4B",   x"2E",   x"81",   x"E4",   x"1C",   x"79",   x"D6",   x"B3", 
  x"E5",   x"80",   x"2F",   x"4A",   x"B2",   x"D7",   x"78",   x"1D", 
  x"D4",   x"B1",   x"1E",   x"7B",   x"83",   x"E6",   x"49",   x"2C", 
  x"7A",   x"1F",   x"B0",   x"D5",   x"2D",   x"48",   x"E7",   x"82", 
  x"B6",   x"D3",   x"7C",   x"19",   x"E1",   x"84",   x"2B",   x"4E", 
  x"18",   x"7D",   x"D2",   x"B7",   x"4F",   x"2A",   x"85",   x"E0", 
  x"29",   x"4C",   x"E3",   x"86",   x"7E",   x"1B",   x"B4",   x"D1", 
  x"87",   x"E2",   x"4D",   x"28",   x"D0",   x"B5",   x"1A",   x"7F", 
  x"00",   x"66",   x"CC",   x"AA",   x"5B",   x"3D",   x"97",   x"F1", 
  x"B6",   x"D0",   x"7A",   x"1C",   x"ED",   x"8B",   x"21",   x"47", 
  x"AF",   x"C9",   x"63",   x"05",   x"F4",   x"92",   x"38",   x"5E", 
  x"19",   x"7F",   x"D5",   x"B3",   x"42",   x"24",   x"8E",   x"E8", 
  x"9D",   x"FB",   x"51",   x"37",   x"C6",   x"A0",   x"0A",   x"6C", 
  x"2B",   x"4D",   x"E7",   x"81",   x"70",   x"16",   x"BC",   x"DA", 
  x"32",   x"54",   x"FE",   x"98",   x"69",   x"0F",   x"A5",   x"C3", 
  x"84",   x"E2",   x"48",   x"2E",   x"DF",   x"B9",   x"13",   x"75", 
  x"F9",   x"9F",   x"35",   x"53",   x"A2",   x"C4",   x"6E",   x"08", 
  x"4F",   x"29",   x"83",   x"E5",   x"14",   x"72",   x"D8",   x"BE", 
  x"56",   x"30",   x"9A",   x"FC",   x"0D",   x"6B",   x"C1",   x"A7", 
  x"E0",   x"86",   x"2C",   x"4A",   x"BB",   x"DD",   x"77",   x"11", 
  x"64",   x"02",   x"A8",   x"CE",   x"3F",   x"59",   x"F3",   x"95", 
  x"D2",   x"B4",   x"1E",   x"78",   x"89",   x"EF",   x"45",   x"23", 
  x"CB",   x"AD",   x"07",   x"61",   x"90",   x"F6",   x"5C",   x"3A", 
  x"7D",   x"1B",   x"B1",   x"D7",   x"26",   x"40",   x"EA",   x"8C", 
  x"31",   x"57",   x"FD",   x"9B",   x"6A",   x"0C",   x"A6",   x"C0", 
  x"87",   x"E1",   x"4B",   x"2D",   x"DC",   x"BA",   x"10",   x"76", 
  x"9E",   x"F8",   x"52",   x"34",   x"C5",   x"A3",   x"09",   x"6F", 
  x"28",   x"4E",   x"E4",   x"82",   x"73",   x"15",   x"BF",   x"D9", 
  x"AC",   x"CA",   x"60",   x"06",   x"F7",   x"91",   x"3B",   x"5D", 
  x"1A",   x"7C",   x"D6",   x"B0",   x"41",   x"27",   x"8D",   x"EB", 
  x"03",   x"65",   x"CF",   x"A9",   x"58",   x"3E",   x"94",   x"F2", 
  x"B5",   x"D3",   x"79",   x"1F",   x"EE",   x"88",   x"22",   x"44", 
  x"C8",   x"AE",   x"04",   x"62",   x"93",   x"F5",   x"5F",   x"39", 
  x"7E",   x"18",   x"B2",   x"D4",   x"25",   x"43",   x"E9",   x"8F", 
  x"67",   x"01",   x"AB",   x"CD",   x"3C",   x"5A",   x"F0",   x"96", 
  x"D1",   x"B7",   x"1D",   x"7B",   x"8A",   x"EC",   x"46",   x"20", 
  x"55",   x"33",   x"99",   x"FF",   x"0E",   x"68",   x"C2",   x"A4", 
  x"E3",   x"85",   x"2F",   x"49",   x"B8",   x"DE",   x"74",   x"12", 
  x"FA",   x"9C",   x"36",   x"50",   x"A1",   x"C7",   x"6D",   x"0B", 
  x"4C",   x"2A",   x"80",   x"E6",   x"17",   x"71",   x"DB",   x"BD", 
  x"00",   x"67",   x"CE",   x"A9",   x"5F",   x"38",   x"91",   x"F6", 
  x"BE",   x"D9",   x"70",   x"17",   x"E1",   x"86",   x"2F",   x"48", 
  x"BF",   x"D8",   x"71",   x"16",   x"E0",   x"87",   x"2E",   x"49", 
  x"01",   x"66",   x"CF",   x"A8",   x"5E",   x"39",   x"90",   x"F7", 
  x"BD",   x"DA",   x"73",   x"14",   x"E2",   x"85",   x"2C",   x"4B", 
  x"03",   x"64",   x"CD",   x"AA",   x"5C",   x"3B",   x"92",   x"F5", 
  x"02",   x"65",   x"CC",   x"AB",   x"5D",   x"3A",   x"93",   x"F4", 
  x"BC",   x"DB",   x"72",   x"15",   x"E3",   x"84",   x"2D",   x"4A", 
  x"B9",   x"DE",   x"77",   x"10",   x"E6",   x"81",   x"28",   x"4F", 
  x"07",   x"60",   x"C9",   x"AE",   x"58",   x"3F",   x"96",   x"F1", 
  x"06",   x"61",   x"C8",   x"AF",   x"59",   x"3E",   x"97",   x"F0", 
  x"B8",   x"DF",   x"76",   x"11",   x"E7",   x"80",   x"29",   x"4E", 
  x"04",   x"63",   x"CA",   x"AD",   x"5B",   x"3C",   x"95",   x"F2", 
  x"BA",   x"DD",   x"74",   x"13",   x"E5",   x"82",   x"2B",   x"4C", 
  x"BB",   x"DC",   x"75",   x"12",   x"E4",   x"83",   x"2A",   x"4D", 
  x"05",   x"62",   x"CB",   x"AC",   x"5A",   x"3D",   x"94",   x"F3", 
  x"B1",   x"D6",   x"7F",   x"18",   x"EE",   x"89",   x"20",   x"47", 
  x"0F",   x"68",   x"C1",   x"A6",   x"50",   x"37",   x"9E",   x"F9", 
  x"0E",   x"69",   x"C0",   x"A7",   x"51",   x"36",   x"9F",   x"F8", 
  x"B0",   x"D7",   x"7E",   x"19",   x"EF",   x"88",   x"21",   x"46", 
  x"0C",   x"6B",   x"C2",   x"A5",   x"53",   x"34",   x"9D",   x"FA", 
  x"B2",   x"D5",   x"7C",   x"1B",   x"ED",   x"8A",   x"23",   x"44", 
  x"B3",   x"D4",   x"7D",   x"1A",   x"EC",   x"8B",   x"22",   x"45", 
  x"0D",   x"6A",   x"C3",   x"A4",   x"52",   x"35",   x"9C",   x"FB", 
  x"08",   x"6F",   x"C6",   x"A1",   x"57",   x"30",   x"99",   x"FE", 
  x"B6",   x"D1",   x"78",   x"1F",   x"E9",   x"8E",   x"27",   x"40", 
  x"B7",   x"D0",   x"79",   x"1E",   x"E8",   x"8F",   x"26",   x"41", 
  x"09",   x"6E",   x"C7",   x"A0",   x"56",   x"31",   x"98",   x"FF", 
  x"B5",   x"D2",   x"7B",   x"1C",   x"EA",   x"8D",   x"24",   x"43", 
  x"0B",   x"6C",   x"C5",   x"A2",   x"54",   x"33",   x"9A",   x"FD", 
  x"0A",   x"6D",   x"C4",   x"A3",   x"55",   x"32",   x"9B",   x"FC", 
  x"B4",   x"D3",   x"7A",   x"1D",   x"EB",   x"8C",   x"25",   x"42", 
  x"00",   x"68",   x"D0",   x"B8",   x"63",   x"0B",   x"B3",   x"DB", 
  x"C6",   x"AE",   x"16",   x"7E",   x"A5",   x"CD",   x"75",   x"1D", 
  x"4F",   x"27",   x"9F",   x"F7",   x"2C",   x"44",   x"FC",   x"94", 
  x"89",   x"E1",   x"59",   x"31",   x"EA",   x"82",   x"3A",   x"52", 
  x"9E",   x"F6",   x"4E",   x"26",   x"FD",   x"95",   x"2D",   x"45", 
  x"58",   x"30",   x"88",   x"E0",   x"3B",   x"53",   x"EB",   x"83", 
  x"D1",   x"B9",   x"01",   x"69",   x"B2",   x"DA",   x"62",   x"0A", 
  x"17",   x"7F",   x"C7",   x"AF",   x"74",   x"1C",   x"A4",   x"CC", 
  x"FF",   x"97",   x"2F",   x"47",   x"9C",   x"F4",   x"4C",   x"24", 
  x"39",   x"51",   x"E9",   x"81",   x"5A",   x"32",   x"8A",   x"E2", 
  x"B0",   x"D8",   x"60",   x"08",   x"D3",   x"BB",   x"03",   x"6B", 
  x"76",   x"1E",   x"A6",   x"CE",   x"15",   x"7D",   x"C5",   x"AD", 
  x"61",   x"09",   x"B1",   x"D9",   x"02",   x"6A",   x"D2",   x"BA", 
  x"A7",   x"CF",   x"77",   x"1F",   x"C4",   x"AC",   x"14",   x"7C", 
  x"2E",   x"46",   x"FE",   x"96",   x"4D",   x"25",   x"9D",   x"F5", 
  x"E8",   x"80",   x"38",   x"50",   x"8B",   x"E3",   x"5B",   x"33", 
  x"3D",   x"55",   x"ED",   x"85",   x"5E",   x"36",   x"8E",   x"E6", 
  x"FB",   x"93",   x"2B",   x"43",   x"98",   x"F0",   x"48",   x"20", 
  x"72",   x"1A",   x"A2",   x"CA",   x"11",   x"79",   x"C1",   x"A9", 
  x"B4",   x"DC",   x"64",   x"0C",   x"D7",   x"BF",   x"07",   x"6F", 
  x"A3",   x"CB",   x"73",   x"1B",   x"C0",   x"A8",   x"10",   x"78", 
  x"65",   x"0D",   x"B5",   x"DD",   x"06",   x"6E",   x"D6",   x"BE", 
  x"EC",   x"84",   x"3C",   x"54",   x"8F",   x"E7",   x"5F",   x"37", 
  x"2A",   x"42",   x"FA",   x"92",   x"49",   x"21",   x"99",   x"F1", 
  x"C2",   x"AA",   x"12",   x"7A",   x"A1",   x"C9",   x"71",   x"19", 
  x"04",   x"6C",   x"D4",   x"BC",   x"67",   x"0F",   x"B7",   x"DF", 
  x"8D",   x"E5",   x"5D",   x"35",   x"EE",   x"86",   x"3E",   x"56", 
  x"4B",   x"23",   x"9B",   x"F3",   x"28",   x"40",   x"F8",   x"90", 
  x"5C",   x"34",   x"8C",   x"E4",   x"3F",   x"57",   x"EF",   x"87", 
  x"9A",   x"F2",   x"4A",   x"22",   x"F9",   x"91",   x"29",   x"41", 
  x"13",   x"7B",   x"C3",   x"AB",   x"70",   x"18",   x"A0",   x"C8", 
  x"D5",   x"BD",   x"05",   x"6D",   x"B6",   x"DE",   x"66",   x"0E", 
  x"00",   x"69",   x"D2",   x"BB",   x"67",   x"0E",   x"B5",   x"DC", 
  x"CE",   x"A7",   x"1C",   x"75",   x"A9",   x"C0",   x"7B",   x"12", 
  x"5F",   x"36",   x"8D",   x"E4",   x"38",   x"51",   x"EA",   x"83", 
  x"91",   x"F8",   x"43",   x"2A",   x"F6",   x"9F",   x"24",   x"4D", 
  x"BE",   x"D7",   x"6C",   x"05",   x"D9",   x"B0",   x"0B",   x"62", 
  x"70",   x"19",   x"A2",   x"CB",   x"17",   x"7E",   x"C5",   x"AC", 
  x"E1",   x"88",   x"33",   x"5A",   x"86",   x"EF",   x"54",   x"3D", 
  x"2F",   x"46",   x"FD",   x"94",   x"48",   x"21",   x"9A",   x"F3", 
  x"BF",   x"D6",   x"6D",   x"04",   x"D8",   x"B1",   x"0A",   x"63", 
  x"71",   x"18",   x"A3",   x"CA",   x"16",   x"7F",   x"C4",   x"AD", 
  x"E0",   x"89",   x"32",   x"5B",   x"87",   x"EE",   x"55",   x"3C", 
  x"2E",   x"47",   x"FC",   x"95",   x"49",   x"20",   x"9B",   x"F2", 
  x"01",   x"68",   x"D3",   x"BA",   x"66",   x"0F",   x"B4",   x"DD", 
  x"CF",   x"A6",   x"1D",   x"74",   x"A8",   x"C1",   x"7A",   x"13", 
  x"5E",   x"37",   x"8C",   x"E5",   x"39",   x"50",   x"EB",   x"82", 
  x"90",   x"F9",   x"42",   x"2B",   x"F7",   x"9E",   x"25",   x"4C", 
  x"BD",   x"D4",   x"6F",   x"06",   x"DA",   x"B3",   x"08",   x"61", 
  x"73",   x"1A",   x"A1",   x"C8",   x"14",   x"7D",   x"C6",   x"AF", 
  x"E2",   x"8B",   x"30",   x"59",   x"85",   x"EC",   x"57",   x"3E", 
  x"2C",   x"45",   x"FE",   x"97",   x"4B",   x"22",   x"99",   x"F0", 
  x"03",   x"6A",   x"D1",   x"B8",   x"64",   x"0D",   x"B6",   x"DF", 
  x"CD",   x"A4",   x"1F",   x"76",   x"AA",   x"C3",   x"78",   x"11", 
  x"5C",   x"35",   x"8E",   x"E7",   x"3B",   x"52",   x"E9",   x"80", 
  x"92",   x"FB",   x"40",   x"29",   x"F5",   x"9C",   x"27",   x"4E", 
  x"02",   x"6B",   x"D0",   x"B9",   x"65",   x"0C",   x"B7",   x"DE", 
  x"CC",   x"A5",   x"1E",   x"77",   x"AB",   x"C2",   x"79",   x"10", 
  x"5D",   x"34",   x"8F",   x"E6",   x"3A",   x"53",   x"E8",   x"81", 
  x"93",   x"FA",   x"41",   x"28",   x"F4",   x"9D",   x"26",   x"4F", 
  x"BC",   x"D5",   x"6E",   x"07",   x"DB",   x"B2",   x"09",   x"60", 
  x"72",   x"1B",   x"A0",   x"C9",   x"15",   x"7C",   x"C7",   x"AE", 
  x"E3",   x"8A",   x"31",   x"58",   x"84",   x"ED",   x"56",   x"3F", 
  x"2D",   x"44",   x"FF",   x"96",   x"4A",   x"23",   x"98",   x"F1", 
  x"00",   x"6A",   x"D4",   x"BE",   x"6B",   x"01",   x"BF",   x"D5", 
  x"D6",   x"BC",   x"02",   x"68",   x"BD",   x"D7",   x"69",   x"03", 
  x"6F",   x"05",   x"BB",   x"D1",   x"04",   x"6E",   x"D0",   x"BA", 
  x"B9",   x"D3",   x"6D",   x"07",   x"D2",   x"B8",   x"06",   x"6C", 
  x"DE",   x"B4",   x"0A",   x"60",   x"B5",   x"DF",   x"61",   x"0B", 
  x"08",   x"62",   x"DC",   x"B6",   x"63",   x"09",   x"B7",   x"DD", 
  x"B1",   x"DB",   x"65",   x"0F",   x"DA",   x"B0",   x"0E",   x"64", 
  x"67",   x"0D",   x"B3",   x"D9",   x"0C",   x"66",   x"D8",   x"B2", 
  x"7F",   x"15",   x"AB",   x"C1",   x"14",   x"7E",   x"C0",   x"AA", 
  x"A9",   x"C3",   x"7D",   x"17",   x"C2",   x"A8",   x"16",   x"7C", 
  x"10",   x"7A",   x"C4",   x"AE",   x"7B",   x"11",   x"AF",   x"C5", 
  x"C6",   x"AC",   x"12",   x"78",   x"AD",   x"C7",   x"79",   x"13", 
  x"A1",   x"CB",   x"75",   x"1F",   x"CA",   x"A0",   x"1E",   x"74", 
  x"77",   x"1D",   x"A3",   x"C9",   x"1C",   x"76",   x"C8",   x"A2", 
  x"CE",   x"A4",   x"1A",   x"70",   x"A5",   x"CF",   x"71",   x"1B", 
  x"18",   x"72",   x"CC",   x"A6",   x"73",   x"19",   x"A7",   x"CD", 
  x"FE",   x"94",   x"2A",   x"40",   x"95",   x"FF",   x"41",   x"2B", 
  x"28",   x"42",   x"FC",   x"96",   x"43",   x"29",   x"97",   x"FD", 
  x"91",   x"FB",   x"45",   x"2F",   x"FA",   x"90",   x"2E",   x"44", 
  x"47",   x"2D",   x"93",   x"F9",   x"2C",   x"46",   x"F8",   x"92", 
  x"20",   x"4A",   x"F4",   x"9E",   x"4B",   x"21",   x"9F",   x"F5", 
  x"F6",   x"9C",   x"22",   x"48",   x"9D",   x"F7",   x"49",   x"23", 
  x"4F",   x"25",   x"9B",   x"F1",   x"24",   x"4E",   x"F0",   x"9A", 
  x"99",   x"F3",   x"4D",   x"27",   x"F2",   x"98",   x"26",   x"4C", 
  x"81",   x"EB",   x"55",   x"3F",   x"EA",   x"80",   x"3E",   x"54", 
  x"57",   x"3D",   x"83",   x"E9",   x"3C",   x"56",   x"E8",   x"82", 
  x"EE",   x"84",   x"3A",   x"50",   x"85",   x"EF",   x"51",   x"3B", 
  x"38",   x"52",   x"EC",   x"86",   x"53",   x"39",   x"87",   x"ED", 
  x"5F",   x"35",   x"8B",   x"E1",   x"34",   x"5E",   x"E0",   x"8A", 
  x"89",   x"E3",   x"5D",   x"37",   x"E2",   x"88",   x"36",   x"5C", 
  x"30",   x"5A",   x"E4",   x"8E",   x"5B",   x"31",   x"8F",   x"E5", 
  x"E6",   x"8C",   x"32",   x"58",   x"8D",   x"E7",   x"59",   x"33", 
  x"00",   x"6B",   x"D6",   x"BD",   x"6F",   x"04",   x"B9",   x"D2", 
  x"DE",   x"B5",   x"08",   x"63",   x"B1",   x"DA",   x"67",   x"0C", 
  x"7F",   x"14",   x"A9",   x"C2",   x"10",   x"7B",   x"C6",   x"AD", 
  x"A1",   x"CA",   x"77",   x"1C",   x"CE",   x"A5",   x"18",   x"73", 
  x"FE",   x"95",   x"28",   x"43",   x"91",   x"FA",   x"47",   x"2C", 
  x"20",   x"4B",   x"F6",   x"9D",   x"4F",   x"24",   x"99",   x"F2", 
  x"81",   x"EA",   x"57",   x"3C",   x"EE",   x"85",   x"38",   x"53", 
  x"5F",   x"34",   x"89",   x"E2",   x"30",   x"5B",   x"E6",   x"8D", 
  x"3F",   x"54",   x"E9",   x"82",   x"50",   x"3B",   x"86",   x"ED", 
  x"E1",   x"8A",   x"37",   x"5C",   x"8E",   x"E5",   x"58",   x"33", 
  x"40",   x"2B",   x"96",   x"FD",   x"2F",   x"44",   x"F9",   x"92", 
  x"9E",   x"F5",   x"48",   x"23",   x"F1",   x"9A",   x"27",   x"4C", 
  x"C1",   x"AA",   x"17",   x"7C",   x"AE",   x"C5",   x"78",   x"13", 
  x"1F",   x"74",   x"C9",   x"A2",   x"70",   x"1B",   x"A6",   x"CD", 
  x"BE",   x"D5",   x"68",   x"03",   x"D1",   x"BA",   x"07",   x"6C", 
  x"60",   x"0B",   x"B6",   x"DD",   x"0F",   x"64",   x"D9",   x"B2", 
  x"7E",   x"15",   x"A8",   x"C3",   x"11",   x"7A",   x"C7",   x"AC", 
  x"A0",   x"CB",   x"76",   x"1D",   x"CF",   x"A4",   x"19",   x"72", 
  x"01",   x"6A",   x"D7",   x"BC",   x"6E",   x"05",   x"B8",   x"D3", 
  x"DF",   x"B4",   x"09",   x"62",   x"B0",   x"DB",   x"66",   x"0D", 
  x"80",   x"EB",   x"56",   x"3D",   x"EF",   x"84",   x"39",   x"52", 
  x"5E",   x"35",   x"88",   x"E3",   x"31",   x"5A",   x"E7",   x"8C", 
  x"FF",   x"94",   x"29",   x"42",   x"90",   x"FB",   x"46",   x"2D", 
  x"21",   x"4A",   x"F7",   x"9C",   x"4E",   x"25",   x"98",   x"F3", 
  x"41",   x"2A",   x"97",   x"FC",   x"2E",   x"45",   x"F8",   x"93", 
  x"9F",   x"F4",   x"49",   x"22",   x"F0",   x"9B",   x"26",   x"4D", 
  x"3E",   x"55",   x"E8",   x"83",   x"51",   x"3A",   x"87",   x"EC", 
  x"E0",   x"8B",   x"36",   x"5D",   x"8F",   x"E4",   x"59",   x"32", 
  x"BF",   x"D4",   x"69",   x"02",   x"D0",   x"BB",   x"06",   x"6D", 
  x"61",   x"0A",   x"B7",   x"DC",   x"0E",   x"65",   x"D8",   x"B3", 
  x"C0",   x"AB",   x"16",   x"7D",   x"AF",   x"C4",   x"79",   x"12", 
  x"1E",   x"75",   x"C8",   x"A3",   x"71",   x"1A",   x"A7",   x"CC", 
  x"00",   x"6C",   x"D8",   x"B4",   x"73",   x"1F",   x"AB",   x"C7", 
  x"E6",   x"8A",   x"3E",   x"52",   x"95",   x"F9",   x"4D",   x"21", 
  x"0F",   x"63",   x"D7",   x"BB",   x"7C",   x"10",   x"A4",   x"C8", 
  x"E9",   x"85",   x"31",   x"5D",   x"9A",   x"F6",   x"42",   x"2E", 
  x"1E",   x"72",   x"C6",   x"AA",   x"6D",   x"01",   x"B5",   x"D9", 
  x"F8",   x"94",   x"20",   x"4C",   x"8B",   x"E7",   x"53",   x"3F", 
  x"11",   x"7D",   x"C9",   x"A5",   x"62",   x"0E",   x"BA",   x"D6", 
  x"F7",   x"9B",   x"2F",   x"43",   x"84",   x"E8",   x"5C",   x"30", 
  x"3C",   x"50",   x"E4",   x"88",   x"4F",   x"23",   x"97",   x"FB", 
  x"DA",   x"B6",   x"02",   x"6E",   x"A9",   x"C5",   x"71",   x"1D", 
  x"33",   x"5F",   x"EB",   x"87",   x"40",   x"2C",   x"98",   x"F4", 
  x"D5",   x"B9",   x"0D",   x"61",   x"A6",   x"CA",   x"7E",   x"12", 
  x"22",   x"4E",   x"FA",   x"96",   x"51",   x"3D",   x"89",   x"E5", 
  x"C4",   x"A8",   x"1C",   x"70",   x"B7",   x"DB",   x"6F",   x"03", 
  x"2D",   x"41",   x"F5",   x"99",   x"5E",   x"32",   x"86",   x"EA", 
  x"CB",   x"A7",   x"13",   x"7F",   x"B8",   x"D4",   x"60",   x"0C", 
  x"78",   x"14",   x"A0",   x"CC",   x"0B",   x"67",   x"D3",   x"BF", 
  x"9E",   x"F2",   x"46",   x"2A",   x"ED",   x"81",   x"35",   x"59", 
  x"77",   x"1B",   x"AF",   x"C3",   x"04",   x"68",   x"DC",   x"B0", 
  x"91",   x"FD",   x"49",   x"25",   x"E2",   x"8E",   x"3A",   x"56", 
  x"66",   x"0A",   x"BE",   x"D2",   x"15",   x"79",   x"CD",   x"A1", 
  x"80",   x"EC",   x"58",   x"34",   x"F3",   x"9F",   x"2B",   x"47", 
  x"69",   x"05",   x"B1",   x"DD",   x"1A",   x"76",   x"C2",   x"AE", 
  x"8F",   x"E3",   x"57",   x"3B",   x"FC",   x"90",   x"24",   x"48", 
  x"44",   x"28",   x"9C",   x"F0",   x"37",   x"5B",   x"EF",   x"83", 
  x"A2",   x"CE",   x"7A",   x"16",   x"D1",   x"BD",   x"09",   x"65", 
  x"4B",   x"27",   x"93",   x"FF",   x"38",   x"54",   x"E0",   x"8C", 
  x"AD",   x"C1",   x"75",   x"19",   x"DE",   x"B2",   x"06",   x"6A", 
  x"5A",   x"36",   x"82",   x"EE",   x"29",   x"45",   x"F1",   x"9D", 
  x"BC",   x"D0",   x"64",   x"08",   x"CF",   x"A3",   x"17",   x"7B", 
  x"55",   x"39",   x"8D",   x"E1",   x"26",   x"4A",   x"FE",   x"92", 
  x"B3",   x"DF",   x"6B",   x"07",   x"C0",   x"AC",   x"18",   x"74", 
  x"00",   x"6D",   x"DA",   x"B7",   x"77",   x"1A",   x"AD",   x"C0", 
  x"EE",   x"83",   x"34",   x"59",   x"99",   x"F4",   x"43",   x"2E", 
  x"1F",   x"72",   x"C5",   x"A8",   x"68",   x"05",   x"B2",   x"DF", 
  x"F1",   x"9C",   x"2B",   x"46",   x"86",   x"EB",   x"5C",   x"31", 
  x"3E",   x"53",   x"E4",   x"89",   x"49",   x"24",   x"93",   x"FE", 
  x"D0",   x"BD",   x"0A",   x"67",   x"A7",   x"CA",   x"7D",   x"10", 
  x"21",   x"4C",   x"FB",   x"96",   x"56",   x"3B",   x"8C",   x"E1", 
  x"CF",   x"A2",   x"15",   x"78",   x"B8",   x"D5",   x"62",   x"0F", 
  x"7C",   x"11",   x"A6",   x"CB",   x"0B",   x"66",   x"D1",   x"BC", 
  x"92",   x"FF",   x"48",   x"25",   x"E5",   x"88",   x"3F",   x"52", 
  x"63",   x"0E",   x"B9",   x"D4",   x"14",   x"79",   x"CE",   x"A3", 
  x"8D",   x"E0",   x"57",   x"3A",   x"FA",   x"97",   x"20",   x"4D", 
  x"42",   x"2F",   x"98",   x"F5",   x"35",   x"58",   x"EF",   x"82", 
  x"AC",   x"C1",   x"76",   x"1B",   x"DB",   x"B6",   x"01",   x"6C", 
  x"5D",   x"30",   x"87",   x"EA",   x"2A",   x"47",   x"F0",   x"9D", 
  x"B3",   x"DE",   x"69",   x"04",   x"C4",   x"A9",   x"1E",   x"73", 
  x"F8",   x"95",   x"22",   x"4F",   x"8F",   x"E2",   x"55",   x"38", 
  x"16",   x"7B",   x"CC",   x"A1",   x"61",   x"0C",   x"BB",   x"D6", 
  x"E7",   x"8A",   x"3D",   x"50",   x"90",   x"FD",   x"4A",   x"27", 
  x"09",   x"64",   x"D3",   x"BE",   x"7E",   x"13",   x"A4",   x"C9", 
  x"C6",   x"AB",   x"1C",   x"71",   x"B1",   x"DC",   x"6B",   x"06", 
  x"28",   x"45",   x"F2",   x"9F",   x"5F",   x"32",   x"85",   x"E8", 
  x"D9",   x"B4",   x"03",   x"6E",   x"AE",   x"C3",   x"74",   x"19", 
  x"37",   x"5A",   x"ED",   x"80",   x"40",   x"2D",   x"9A",   x"F7", 
  x"84",   x"E9",   x"5E",   x"33",   x"F3",   x"9E",   x"29",   x"44", 
  x"6A",   x"07",   x"B0",   x"DD",   x"1D",   x"70",   x"C7",   x"AA", 
  x"9B",   x"F6",   x"41",   x"2C",   x"EC",   x"81",   x"36",   x"5B", 
  x"75",   x"18",   x"AF",   x"C2",   x"02",   x"6F",   x"D8",   x"B5", 
  x"BA",   x"D7",   x"60",   x"0D",   x"CD",   x"A0",   x"17",   x"7A", 
  x"54",   x"39",   x"8E",   x"E3",   x"23",   x"4E",   x"F9",   x"94", 
  x"A5",   x"C8",   x"7F",   x"12",   x"D2",   x"BF",   x"08",   x"65", 
  x"4B",   x"26",   x"91",   x"FC",   x"3C",   x"51",   x"E6",   x"8B", 
  x"00",   x"6E",   x"DC",   x"B2",   x"7B",   x"15",   x"A7",   x"C9", 
  x"F6",   x"98",   x"2A",   x"44",   x"8D",   x"E3",   x"51",   x"3F", 
  x"2F",   x"41",   x"F3",   x"9D",   x"54",   x"3A",   x"88",   x"E6", 
  x"D9",   x"B7",   x"05",   x"6B",   x"A2",   x"CC",   x"7E",   x"10", 
  x"5E",   x"30",   x"82",   x"EC",   x"25",   x"4B",   x"F9",   x"97", 
  x"A8",   x"C6",   x"74",   x"1A",   x"D3",   x"BD",   x"0F",   x"61", 
  x"71",   x"1F",   x"AD",   x"C3",   x"0A",   x"64",   x"D6",   x"B8", 
  x"87",   x"E9",   x"5B",   x"35",   x"FC",   x"92",   x"20",   x"4E", 
  x"BC",   x"D2",   x"60",   x"0E",   x"C7",   x"A9",   x"1B",   x"75", 
  x"4A",   x"24",   x"96",   x"F8",   x"31",   x"5F",   x"ED",   x"83", 
  x"93",   x"FD",   x"4F",   x"21",   x"E8",   x"86",   x"34",   x"5A", 
  x"65",   x"0B",   x"B9",   x"D7",   x"1E",   x"70",   x"C2",   x"AC", 
  x"E2",   x"8C",   x"3E",   x"50",   x"99",   x"F7",   x"45",   x"2B", 
  x"14",   x"7A",   x"C8",   x"A6",   x"6F",   x"01",   x"B3",   x"DD", 
  x"CD",   x"A3",   x"11",   x"7F",   x"B6",   x"D8",   x"6A",   x"04", 
  x"3B",   x"55",   x"E7",   x"89",   x"40",   x"2E",   x"9C",   x"F2", 
  x"BB",   x"D5",   x"67",   x"09",   x"C0",   x"AE",   x"1C",   x"72", 
  x"4D",   x"23",   x"91",   x"FF",   x"36",   x"58",   x"EA",   x"84", 
  x"94",   x"FA",   x"48",   x"26",   x"EF",   x"81",   x"33",   x"5D", 
  x"62",   x"0C",   x"BE",   x"D0",   x"19",   x"77",   x"C5",   x"AB", 
  x"E5",   x"8B",   x"39",   x"57",   x"9E",   x"F0",   x"42",   x"2C", 
  x"13",   x"7D",   x"CF",   x"A1",   x"68",   x"06",   x"B4",   x"DA", 
  x"CA",   x"A4",   x"16",   x"78",   x"B1",   x"DF",   x"6D",   x"03", 
  x"3C",   x"52",   x"E0",   x"8E",   x"47",   x"29",   x"9B",   x"F5", 
  x"07",   x"69",   x"DB",   x"B5",   x"7C",   x"12",   x"A0",   x"CE", 
  x"F1",   x"9F",   x"2D",   x"43",   x"8A",   x"E4",   x"56",   x"38", 
  x"28",   x"46",   x"F4",   x"9A",   x"53",   x"3D",   x"8F",   x"E1", 
  x"DE",   x"B0",   x"02",   x"6C",   x"A5",   x"CB",   x"79",   x"17", 
  x"59",   x"37",   x"85",   x"EB",   x"22",   x"4C",   x"FE",   x"90", 
  x"AF",   x"C1",   x"73",   x"1D",   x"D4",   x"BA",   x"08",   x"66", 
  x"76",   x"18",   x"AA",   x"C4",   x"0D",   x"63",   x"D1",   x"BF", 
  x"80",   x"EE",   x"5C",   x"32",   x"FB",   x"95",   x"27",   x"49", 
  x"00",   x"6F",   x"DE",   x"B1",   x"7F",   x"10",   x"A1",   x"CE", 
  x"FE",   x"91",   x"20",   x"4F",   x"81",   x"EE",   x"5F",   x"30", 
  x"3F",   x"50",   x"E1",   x"8E",   x"40",   x"2F",   x"9E",   x"F1", 
  x"C1",   x"AE",   x"1F",   x"70",   x"BE",   x"D1",   x"60",   x"0F", 
  x"7E",   x"11",   x"A0",   x"CF",   x"01",   x"6E",   x"DF",   x"B0", 
  x"80",   x"EF",   x"5E",   x"31",   x"FF",   x"90",   x"21",   x"4E", 
  x"41",   x"2E",   x"9F",   x"F0",   x"3E",   x"51",   x"E0",   x"8F", 
  x"BF",   x"D0",   x"61",   x"0E",   x"C0",   x"AF",   x"1E",   x"71", 
  x"FC",   x"93",   x"22",   x"4D",   x"83",   x"EC",   x"5D",   x"32", 
  x"02",   x"6D",   x"DC",   x"B3",   x"7D",   x"12",   x"A3",   x"CC", 
  x"C3",   x"AC",   x"1D",   x"72",   x"BC",   x"D3",   x"62",   x"0D", 
  x"3D",   x"52",   x"E3",   x"8C",   x"42",   x"2D",   x"9C",   x"F3", 
  x"82",   x"ED",   x"5C",   x"33",   x"FD",   x"92",   x"23",   x"4C", 
  x"7C",   x"13",   x"A2",   x"CD",   x"03",   x"6C",   x"DD",   x"B2", 
  x"BD",   x"D2",   x"63",   x"0C",   x"C2",   x"AD",   x"1C",   x"73", 
  x"43",   x"2C",   x"9D",   x"F2",   x"3C",   x"53",   x"E2",   x"8D", 
  x"3B",   x"54",   x"E5",   x"8A",   x"44",   x"2B",   x"9A",   x"F5", 
  x"C5",   x"AA",   x"1B",   x"74",   x"BA",   x"D5",   x"64",   x"0B", 
  x"04",   x"6B",   x"DA",   x"B5",   x"7B",   x"14",   x"A5",   x"CA", 
  x"FA",   x"95",   x"24",   x"4B",   x"85",   x"EA",   x"5B",   x"34", 
  x"45",   x"2A",   x"9B",   x"F4",   x"3A",   x"55",   x"E4",   x"8B", 
  x"BB",   x"D4",   x"65",   x"0A",   x"C4",   x"AB",   x"1A",   x"75", 
  x"7A",   x"15",   x"A4",   x"CB",   x"05",   x"6A",   x"DB",   x"B4", 
  x"84",   x"EB",   x"5A",   x"35",   x"FB",   x"94",   x"25",   x"4A", 
  x"C7",   x"A8",   x"19",   x"76",   x"B8",   x"D7",   x"66",   x"09", 
  x"39",   x"56",   x"E7",   x"88",   x"46",   x"29",   x"98",   x"F7", 
  x"F8",   x"97",   x"26",   x"49",   x"87",   x"E8",   x"59",   x"36", 
  x"06",   x"69",   x"D8",   x"B7",   x"79",   x"16",   x"A7",   x"C8", 
  x"B9",   x"D6",   x"67",   x"08",   x"C6",   x"A9",   x"18",   x"77", 
  x"47",   x"28",   x"99",   x"F6",   x"38",   x"57",   x"E6",   x"89", 
  x"86",   x"E9",   x"58",   x"37",   x"F9",   x"96",   x"27",   x"48", 
  x"78",   x"17",   x"A6",   x"C9",   x"07",   x"68",   x"D9",   x"B6", 
  x"00",   x"70",   x"E0",   x"90",   x"03",   x"73",   x"E3",   x"93", 
  x"06",   x"76",   x"E6",   x"96",   x"05",   x"75",   x"E5",   x"95", 
  x"0C",   x"7C",   x"EC",   x"9C",   x"0F",   x"7F",   x"EF",   x"9F", 
  x"0A",   x"7A",   x"EA",   x"9A",   x"09",   x"79",   x"E9",   x"99", 
  x"18",   x"68",   x"F8",   x"88",   x"1B",   x"6B",   x"FB",   x"8B", 
  x"1E",   x"6E",   x"FE",   x"8E",   x"1D",   x"6D",   x"FD",   x"8D", 
  x"14",   x"64",   x"F4",   x"84",   x"17",   x"67",   x"F7",   x"87", 
  x"12",   x"62",   x"F2",   x"82",   x"11",   x"61",   x"F1",   x"81", 
  x"30",   x"40",   x"D0",   x"A0",   x"33",   x"43",   x"D3",   x"A3", 
  x"36",   x"46",   x"D6",   x"A6",   x"35",   x"45",   x"D5",   x"A5", 
  x"3C",   x"4C",   x"DC",   x"AC",   x"3F",   x"4F",   x"DF",   x"AF", 
  x"3A",   x"4A",   x"DA",   x"AA",   x"39",   x"49",   x"D9",   x"A9", 
  x"28",   x"58",   x"C8",   x"B8",   x"2B",   x"5B",   x"CB",   x"BB", 
  x"2E",   x"5E",   x"CE",   x"BE",   x"2D",   x"5D",   x"CD",   x"BD", 
  x"24",   x"54",   x"C4",   x"B4",   x"27",   x"57",   x"C7",   x"B7", 
  x"22",   x"52",   x"C2",   x"B2",   x"21",   x"51",   x"C1",   x"B1", 
  x"60",   x"10",   x"80",   x"F0",   x"63",   x"13",   x"83",   x"F3", 
  x"66",   x"16",   x"86",   x"F6",   x"65",   x"15",   x"85",   x"F5", 
  x"6C",   x"1C",   x"8C",   x"FC",   x"6F",   x"1F",   x"8F",   x"FF", 
  x"6A",   x"1A",   x"8A",   x"FA",   x"69",   x"19",   x"89",   x"F9", 
  x"78",   x"08",   x"98",   x"E8",   x"7B",   x"0B",   x"9B",   x"EB", 
  x"7E",   x"0E",   x"9E",   x"EE",   x"7D",   x"0D",   x"9D",   x"ED", 
  x"74",   x"04",   x"94",   x"E4",   x"77",   x"07",   x"97",   x"E7", 
  x"72",   x"02",   x"92",   x"E2",   x"71",   x"01",   x"91",   x"E1", 
  x"50",   x"20",   x"B0",   x"C0",   x"53",   x"23",   x"B3",   x"C3", 
  x"56",   x"26",   x"B6",   x"C6",   x"55",   x"25",   x"B5",   x"C5", 
  x"5C",   x"2C",   x"BC",   x"CC",   x"5F",   x"2F",   x"BF",   x"CF", 
  x"5A",   x"2A",   x"BA",   x"CA",   x"59",   x"29",   x"B9",   x"C9", 
  x"48",   x"38",   x"A8",   x"D8",   x"4B",   x"3B",   x"AB",   x"DB", 
  x"4E",   x"3E",   x"AE",   x"DE",   x"4D",   x"3D",   x"AD",   x"DD", 
  x"44",   x"34",   x"A4",   x"D4",   x"47",   x"37",   x"A7",   x"D7", 
  x"42",   x"32",   x"A2",   x"D2",   x"41",   x"31",   x"A1",   x"D1", 
  x"00",   x"71",   x"E2",   x"93",   x"07",   x"76",   x"E5",   x"94", 
  x"0E",   x"7F",   x"EC",   x"9D",   x"09",   x"78",   x"EB",   x"9A", 
  x"1C",   x"6D",   x"FE",   x"8F",   x"1B",   x"6A",   x"F9",   x"88", 
  x"12",   x"63",   x"F0",   x"81",   x"15",   x"64",   x"F7",   x"86", 
  x"38",   x"49",   x"DA",   x"AB",   x"3F",   x"4E",   x"DD",   x"AC", 
  x"36",   x"47",   x"D4",   x"A5",   x"31",   x"40",   x"D3",   x"A2", 
  x"24",   x"55",   x"C6",   x"B7",   x"23",   x"52",   x"C1",   x"B0", 
  x"2A",   x"5B",   x"C8",   x"B9",   x"2D",   x"5C",   x"CF",   x"BE", 
  x"70",   x"01",   x"92",   x"E3",   x"77",   x"06",   x"95",   x"E4", 
  x"7E",   x"0F",   x"9C",   x"ED",   x"79",   x"08",   x"9B",   x"EA", 
  x"6C",   x"1D",   x"8E",   x"FF",   x"6B",   x"1A",   x"89",   x"F8", 
  x"62",   x"13",   x"80",   x"F1",   x"65",   x"14",   x"87",   x"F6", 
  x"48",   x"39",   x"AA",   x"DB",   x"4F",   x"3E",   x"AD",   x"DC", 
  x"46",   x"37",   x"A4",   x"D5",   x"41",   x"30",   x"A3",   x"D2", 
  x"54",   x"25",   x"B6",   x"C7",   x"53",   x"22",   x"B1",   x"C0", 
  x"5A",   x"2B",   x"B8",   x"C9",   x"5D",   x"2C",   x"BF",   x"CE", 
  x"E0",   x"91",   x"02",   x"73",   x"E7",   x"96",   x"05",   x"74", 
  x"EE",   x"9F",   x"0C",   x"7D",   x"E9",   x"98",   x"0B",   x"7A", 
  x"FC",   x"8D",   x"1E",   x"6F",   x"FB",   x"8A",   x"19",   x"68", 
  x"F2",   x"83",   x"10",   x"61",   x"F5",   x"84",   x"17",   x"66", 
  x"D8",   x"A9",   x"3A",   x"4B",   x"DF",   x"AE",   x"3D",   x"4C", 
  x"D6",   x"A7",   x"34",   x"45",   x"D1",   x"A0",   x"33",   x"42", 
  x"C4",   x"B5",   x"26",   x"57",   x"C3",   x"B2",   x"21",   x"50", 
  x"CA",   x"BB",   x"28",   x"59",   x"CD",   x"BC",   x"2F",   x"5E", 
  x"90",   x"E1",   x"72",   x"03",   x"97",   x"E6",   x"75",   x"04", 
  x"9E",   x"EF",   x"7C",   x"0D",   x"99",   x"E8",   x"7B",   x"0A", 
  x"8C",   x"FD",   x"6E",   x"1F",   x"8B",   x"FA",   x"69",   x"18", 
  x"82",   x"F3",   x"60",   x"11",   x"85",   x"F4",   x"67",   x"16", 
  x"A8",   x"D9",   x"4A",   x"3B",   x"AF",   x"DE",   x"4D",   x"3C", 
  x"A6",   x"D7",   x"44",   x"35",   x"A1",   x"D0",   x"43",   x"32", 
  x"B4",   x"C5",   x"56",   x"27",   x"B3",   x"C2",   x"51",   x"20", 
  x"BA",   x"CB",   x"58",   x"29",   x"BD",   x"CC",   x"5F",   x"2E", 
  x"00",   x"72",   x"E4",   x"96",   x"0B",   x"79",   x"EF",   x"9D", 
  x"16",   x"64",   x"F2",   x"80",   x"1D",   x"6F",   x"F9",   x"8B", 
  x"2C",   x"5E",   x"C8",   x"BA",   x"27",   x"55",   x"C3",   x"B1", 
  x"3A",   x"48",   x"DE",   x"AC",   x"31",   x"43",   x"D5",   x"A7", 
  x"58",   x"2A",   x"BC",   x"CE",   x"53",   x"21",   x"B7",   x"C5", 
  x"4E",   x"3C",   x"AA",   x"D8",   x"45",   x"37",   x"A1",   x"D3", 
  x"74",   x"06",   x"90",   x"E2",   x"7F",   x"0D",   x"9B",   x"E9", 
  x"62",   x"10",   x"86",   x"F4",   x"69",   x"1B",   x"8D",   x"FF", 
  x"B0",   x"C2",   x"54",   x"26",   x"BB",   x"C9",   x"5F",   x"2D", 
  x"A6",   x"D4",   x"42",   x"30",   x"AD",   x"DF",   x"49",   x"3B", 
  x"9C",   x"EE",   x"78",   x"0A",   x"97",   x"E5",   x"73",   x"01", 
  x"8A",   x"F8",   x"6E",   x"1C",   x"81",   x"F3",   x"65",   x"17", 
  x"E8",   x"9A",   x"0C",   x"7E",   x"E3",   x"91",   x"07",   x"75", 
  x"FE",   x"8C",   x"1A",   x"68",   x"F5",   x"87",   x"11",   x"63", 
  x"C4",   x"B6",   x"20",   x"52",   x"CF",   x"BD",   x"2B",   x"59", 
  x"D2",   x"A0",   x"36",   x"44",   x"D9",   x"AB",   x"3D",   x"4F", 
  x"A3",   x"D1",   x"47",   x"35",   x"A8",   x"DA",   x"4C",   x"3E", 
  x"B5",   x"C7",   x"51",   x"23",   x"BE",   x"CC",   x"5A",   x"28", 
  x"8F",   x"FD",   x"6B",   x"19",   x"84",   x"F6",   x"60",   x"12", 
  x"99",   x"EB",   x"7D",   x"0F",   x"92",   x"E0",   x"76",   x"04", 
  x"FB",   x"89",   x"1F",   x"6D",   x"F0",   x"82",   x"14",   x"66", 
  x"ED",   x"9F",   x"09",   x"7B",   x"E6",   x"94",   x"02",   x"70", 
  x"D7",   x"A5",   x"33",   x"41",   x"DC",   x"AE",   x"38",   x"4A", 
  x"C1",   x"B3",   x"25",   x"57",   x"CA",   x"B8",   x"2E",   x"5C", 
  x"13",   x"61",   x"F7",   x"85",   x"18",   x"6A",   x"FC",   x"8E", 
  x"05",   x"77",   x"E1",   x"93",   x"0E",   x"7C",   x"EA",   x"98", 
  x"3F",   x"4D",   x"DB",   x"A9",   x"34",   x"46",   x"D0",   x"A2", 
  x"29",   x"5B",   x"CD",   x"BF",   x"22",   x"50",   x"C6",   x"B4", 
  x"4B",   x"39",   x"AF",   x"DD",   x"40",   x"32",   x"A4",   x"D6", 
  x"5D",   x"2F",   x"B9",   x"CB",   x"56",   x"24",   x"B2",   x"C0", 
  x"67",   x"15",   x"83",   x"F1",   x"6C",   x"1E",   x"88",   x"FA", 
  x"71",   x"03",   x"95",   x"E7",   x"7A",   x"08",   x"9E",   x"EC", 
  x"00",   x"73",   x"E6",   x"95",   x"0F",   x"7C",   x"E9",   x"9A", 
  x"1E",   x"6D",   x"F8",   x"8B",   x"11",   x"62",   x"F7",   x"84", 
  x"3C",   x"4F",   x"DA",   x"A9",   x"33",   x"40",   x"D5",   x"A6", 
  x"22",   x"51",   x"C4",   x"B7",   x"2D",   x"5E",   x"CB",   x"B8", 
  x"78",   x"0B",   x"9E",   x"ED",   x"77",   x"04",   x"91",   x"E2", 
  x"66",   x"15",   x"80",   x"F3",   x"69",   x"1A",   x"8F",   x"FC", 
  x"44",   x"37",   x"A2",   x"D1",   x"4B",   x"38",   x"AD",   x"DE", 
  x"5A",   x"29",   x"BC",   x"CF",   x"55",   x"26",   x"B3",   x"C0", 
  x"F0",   x"83",   x"16",   x"65",   x"FF",   x"8C",   x"19",   x"6A", 
  x"EE",   x"9D",   x"08",   x"7B",   x"E1",   x"92",   x"07",   x"74", 
  x"CC",   x"BF",   x"2A",   x"59",   x"C3",   x"B0",   x"25",   x"56", 
  x"D2",   x"A1",   x"34",   x"47",   x"DD",   x"AE",   x"3B",   x"48", 
  x"88",   x"FB",   x"6E",   x"1D",   x"87",   x"F4",   x"61",   x"12", 
  x"96",   x"E5",   x"70",   x"03",   x"99",   x"EA",   x"7F",   x"0C", 
  x"B4",   x"C7",   x"52",   x"21",   x"BB",   x"C8",   x"5D",   x"2E", 
  x"AA",   x"D9",   x"4C",   x"3F",   x"A5",   x"D6",   x"43",   x"30", 
  x"23",   x"50",   x"C5",   x"B6",   x"2C",   x"5F",   x"CA",   x"B9", 
  x"3D",   x"4E",   x"DB",   x"A8",   x"32",   x"41",   x"D4",   x"A7", 
  x"1F",   x"6C",   x"F9",   x"8A",   x"10",   x"63",   x"F6",   x"85", 
  x"01",   x"72",   x"E7",   x"94",   x"0E",   x"7D",   x"E8",   x"9B", 
  x"5B",   x"28",   x"BD",   x"CE",   x"54",   x"27",   x"B2",   x"C1", 
  x"45",   x"36",   x"A3",   x"D0",   x"4A",   x"39",   x"AC",   x"DF", 
  x"67",   x"14",   x"81",   x"F2",   x"68",   x"1B",   x"8E",   x"FD", 
  x"79",   x"0A",   x"9F",   x"EC",   x"76",   x"05",   x"90",   x"E3", 
  x"D3",   x"A0",   x"35",   x"46",   x"DC",   x"AF",   x"3A",   x"49", 
  x"CD",   x"BE",   x"2B",   x"58",   x"C2",   x"B1",   x"24",   x"57", 
  x"EF",   x"9C",   x"09",   x"7A",   x"E0",   x"93",   x"06",   x"75", 
  x"F1",   x"82",   x"17",   x"64",   x"FE",   x"8D",   x"18",   x"6B", 
  x"AB",   x"D8",   x"4D",   x"3E",   x"A4",   x"D7",   x"42",   x"31", 
  x"B5",   x"C6",   x"53",   x"20",   x"BA",   x"C9",   x"5C",   x"2F", 
  x"97",   x"E4",   x"71",   x"02",   x"98",   x"EB",   x"7E",   x"0D", 
  x"89",   x"FA",   x"6F",   x"1C",   x"86",   x"F5",   x"60",   x"13", 
  x"00",   x"74",   x"E8",   x"9C",   x"13",   x"67",   x"FB",   x"8F", 
  x"26",   x"52",   x"CE",   x"BA",   x"35",   x"41",   x"DD",   x"A9", 
  x"4C",   x"38",   x"A4",   x"D0",   x"5F",   x"2B",   x"B7",   x"C3", 
  x"6A",   x"1E",   x"82",   x"F6",   x"79",   x"0D",   x"91",   x"E5", 
  x"98",   x"EC",   x"70",   x"04",   x"8B",   x"FF",   x"63",   x"17", 
  x"BE",   x"CA",   x"56",   x"22",   x"AD",   x"D9",   x"45",   x"31", 
  x"D4",   x"A0",   x"3C",   x"48",   x"C7",   x"B3",   x"2F",   x"5B", 
  x"F2",   x"86",   x"1A",   x"6E",   x"E1",   x"95",   x"09",   x"7D", 
  x"F3",   x"87",   x"1B",   x"6F",   x"E0",   x"94",   x"08",   x"7C", 
  x"D5",   x"A1",   x"3D",   x"49",   x"C6",   x"B2",   x"2E",   x"5A", 
  x"BF",   x"CB",   x"57",   x"23",   x"AC",   x"D8",   x"44",   x"30", 
  x"99",   x"ED",   x"71",   x"05",   x"8A",   x"FE",   x"62",   x"16", 
  x"6B",   x"1F",   x"83",   x"F7",   x"78",   x"0C",   x"90",   x"E4", 
  x"4D",   x"39",   x"A5",   x"D1",   x"5E",   x"2A",   x"B6",   x"C2", 
  x"27",   x"53",   x"CF",   x"BB",   x"34",   x"40",   x"DC",   x"A8", 
  x"01",   x"75",   x"E9",   x"9D",   x"12",   x"66",   x"FA",   x"8E", 
  x"25",   x"51",   x"CD",   x"B9",   x"36",   x"42",   x"DE",   x"AA", 
  x"03",   x"77",   x"EB",   x"9F",   x"10",   x"64",   x"F8",   x"8C", 
  x"69",   x"1D",   x"81",   x"F5",   x"7A",   x"0E",   x"92",   x"E6", 
  x"4F",   x"3B",   x"A7",   x"D3",   x"5C",   x"28",   x"B4",   x"C0", 
  x"BD",   x"C9",   x"55",   x"21",   x"AE",   x"DA",   x"46",   x"32", 
  x"9B",   x"EF",   x"73",   x"07",   x"88",   x"FC",   x"60",   x"14", 
  x"F1",   x"85",   x"19",   x"6D",   x"E2",   x"96",   x"0A",   x"7E", 
  x"D7",   x"A3",   x"3F",   x"4B",   x"C4",   x"B0",   x"2C",   x"58", 
  x"D6",   x"A2",   x"3E",   x"4A",   x"C5",   x"B1",   x"2D",   x"59", 
  x"F0",   x"84",   x"18",   x"6C",   x"E3",   x"97",   x"0B",   x"7F", 
  x"9A",   x"EE",   x"72",   x"06",   x"89",   x"FD",   x"61",   x"15", 
  x"BC",   x"C8",   x"54",   x"20",   x"AF",   x"DB",   x"47",   x"33", 
  x"4E",   x"3A",   x"A6",   x"D2",   x"5D",   x"29",   x"B5",   x"C1", 
  x"68",   x"1C",   x"80",   x"F4",   x"7B",   x"0F",   x"93",   x"E7", 
  x"02",   x"76",   x"EA",   x"9E",   x"11",   x"65",   x"F9",   x"8D", 
  x"24",   x"50",   x"CC",   x"B8",   x"37",   x"43",   x"DF",   x"AB", 
  x"00",   x"75",   x"EA",   x"9F",   x"17",   x"62",   x"FD",   x"88", 
  x"2E",   x"5B",   x"C4",   x"B1",   x"39",   x"4C",   x"D3",   x"A6", 
  x"5C",   x"29",   x"B6",   x"C3",   x"4B",   x"3E",   x"A1",   x"D4", 
  x"72",   x"07",   x"98",   x"ED",   x"65",   x"10",   x"8F",   x"FA", 
  x"B8",   x"CD",   x"52",   x"27",   x"AF",   x"DA",   x"45",   x"30", 
  x"96",   x"E3",   x"7C",   x"09",   x"81",   x"F4",   x"6B",   x"1E", 
  x"E4",   x"91",   x"0E",   x"7B",   x"F3",   x"86",   x"19",   x"6C", 
  x"CA",   x"BF",   x"20",   x"55",   x"DD",   x"A8",   x"37",   x"42", 
  x"B3",   x"C6",   x"59",   x"2C",   x"A4",   x"D1",   x"4E",   x"3B", 
  x"9D",   x"E8",   x"77",   x"02",   x"8A",   x"FF",   x"60",   x"15", 
  x"EF",   x"9A",   x"05",   x"70",   x"F8",   x"8D",   x"12",   x"67", 
  x"C1",   x"B4",   x"2B",   x"5E",   x"D6",   x"A3",   x"3C",   x"49", 
  x"0B",   x"7E",   x"E1",   x"94",   x"1C",   x"69",   x"F6",   x"83", 
  x"25",   x"50",   x"CF",   x"BA",   x"32",   x"47",   x"D8",   x"AD", 
  x"57",   x"22",   x"BD",   x"C8",   x"40",   x"35",   x"AA",   x"DF", 
  x"79",   x"0C",   x"93",   x"E6",   x"6E",   x"1B",   x"84",   x"F1", 
  x"A5",   x"D0",   x"4F",   x"3A",   x"B2",   x"C7",   x"58",   x"2D", 
  x"8B",   x"FE",   x"61",   x"14",   x"9C",   x"E9",   x"76",   x"03", 
  x"F9",   x"8C",   x"13",   x"66",   x"EE",   x"9B",   x"04",   x"71", 
  x"D7",   x"A2",   x"3D",   x"48",   x"C0",   x"B5",   x"2A",   x"5F", 
  x"1D",   x"68",   x"F7",   x"82",   x"0A",   x"7F",   x"E0",   x"95", 
  x"33",   x"46",   x"D9",   x"AC",   x"24",   x"51",   x"CE",   x"BB", 
  x"41",   x"34",   x"AB",   x"DE",   x"56",   x"23",   x"BC",   x"C9", 
  x"6F",   x"1A",   x"85",   x"F0",   x"78",   x"0D",   x"92",   x"E7", 
  x"16",   x"63",   x"FC",   x"89",   x"01",   x"74",   x"EB",   x"9E", 
  x"38",   x"4D",   x"D2",   x"A7",   x"2F",   x"5A",   x"C5",   x"B0", 
  x"4A",   x"3F",   x"A0",   x"D5",   x"5D",   x"28",   x"B7",   x"C2", 
  x"64",   x"11",   x"8E",   x"FB",   x"73",   x"06",   x"99",   x"EC", 
  x"AE",   x"DB",   x"44",   x"31",   x"B9",   x"CC",   x"53",   x"26", 
  x"80",   x"F5",   x"6A",   x"1F",   x"97",   x"E2",   x"7D",   x"08", 
  x"F2",   x"87",   x"18",   x"6D",   x"E5",   x"90",   x"0F",   x"7A", 
  x"DC",   x"A9",   x"36",   x"43",   x"CB",   x"BE",   x"21",   x"54", 
  x"00",   x"76",   x"EC",   x"9A",   x"1B",   x"6D",   x"F7",   x"81", 
  x"36",   x"40",   x"DA",   x"AC",   x"2D",   x"5B",   x"C1",   x"B7", 
  x"6C",   x"1A",   x"80",   x"F6",   x"77",   x"01",   x"9B",   x"ED", 
  x"5A",   x"2C",   x"B6",   x"C0",   x"41",   x"37",   x"AD",   x"DB", 
  x"D8",   x"AE",   x"34",   x"42",   x"C3",   x"B5",   x"2F",   x"59", 
  x"EE",   x"98",   x"02",   x"74",   x"F5",   x"83",   x"19",   x"6F", 
  x"B4",   x"C2",   x"58",   x"2E",   x"AF",   x"D9",   x"43",   x"35", 
  x"82",   x"F4",   x"6E",   x"18",   x"99",   x"EF",   x"75",   x"03", 
  x"73",   x"05",   x"9F",   x"E9",   x"68",   x"1E",   x"84",   x"F2", 
  x"45",   x"33",   x"A9",   x"DF",   x"5E",   x"28",   x"B2",   x"C4", 
  x"1F",   x"69",   x"F3",   x"85",   x"04",   x"72",   x"E8",   x"9E", 
  x"29",   x"5F",   x"C5",   x"B3",   x"32",   x"44",   x"DE",   x"A8", 
  x"AB",   x"DD",   x"47",   x"31",   x"B0",   x"C6",   x"5C",   x"2A", 
  x"9D",   x"EB",   x"71",   x"07",   x"86",   x"F0",   x"6A",   x"1C", 
  x"C7",   x"B1",   x"2B",   x"5D",   x"DC",   x"AA",   x"30",   x"46", 
  x"F1",   x"87",   x"1D",   x"6B",   x"EA",   x"9C",   x"06",   x"70", 
  x"E6",   x"90",   x"0A",   x"7C",   x"FD",   x"8B",   x"11",   x"67", 
  x"D0",   x"A6",   x"3C",   x"4A",   x"CB",   x"BD",   x"27",   x"51", 
  x"8A",   x"FC",   x"66",   x"10",   x"91",   x"E7",   x"7D",   x"0B", 
  x"BC",   x"CA",   x"50",   x"26",   x"A7",   x"D1",   x"4B",   x"3D", 
  x"3E",   x"48",   x"D2",   x"A4",   x"25",   x"53",   x"C9",   x"BF", 
  x"08",   x"7E",   x"E4",   x"92",   x"13",   x"65",   x"FF",   x"89", 
  x"52",   x"24",   x"BE",   x"C8",   x"49",   x"3F",   x"A5",   x"D3", 
  x"64",   x"12",   x"88",   x"FE",   x"7F",   x"09",   x"93",   x"E5", 
  x"95",   x"E3",   x"79",   x"0F",   x"8E",   x"F8",   x"62",   x"14", 
  x"A3",   x"D5",   x"4F",   x"39",   x"B8",   x"CE",   x"54",   x"22", 
  x"F9",   x"8F",   x"15",   x"63",   x"E2",   x"94",   x"0E",   x"78", 
  x"CF",   x"B9",   x"23",   x"55",   x"D4",   x"A2",   x"38",   x"4E", 
  x"4D",   x"3B",   x"A1",   x"D7",   x"56",   x"20",   x"BA",   x"CC", 
  x"7B",   x"0D",   x"97",   x"E1",   x"60",   x"16",   x"8C",   x"FA", 
  x"21",   x"57",   x"CD",   x"BB",   x"3A",   x"4C",   x"D6",   x"A0", 
  x"17",   x"61",   x"FB",   x"8D",   x"0C",   x"7A",   x"E0",   x"96", 
  x"00",   x"77",   x"EE",   x"99",   x"1F",   x"68",   x"F1",   x"86", 
  x"3E",   x"49",   x"D0",   x"A7",   x"21",   x"56",   x"CF",   x"B8", 
  x"7C",   x"0B",   x"92",   x"E5",   x"63",   x"14",   x"8D",   x"FA", 
  x"42",   x"35",   x"AC",   x"DB",   x"5D",   x"2A",   x"B3",   x"C4", 
  x"F8",   x"8F",   x"16",   x"61",   x"E7",   x"90",   x"09",   x"7E", 
  x"C6",   x"B1",   x"28",   x"5F",   x"D9",   x"AE",   x"37",   x"40", 
  x"84",   x"F3",   x"6A",   x"1D",   x"9B",   x"EC",   x"75",   x"02", 
  x"BA",   x"CD",   x"54",   x"23",   x"A5",   x"D2",   x"4B",   x"3C", 
  x"33",   x"44",   x"DD",   x"AA",   x"2C",   x"5B",   x"C2",   x"B5", 
  x"0D",   x"7A",   x"E3",   x"94",   x"12",   x"65",   x"FC",   x"8B", 
  x"4F",   x"38",   x"A1",   x"D6",   x"50",   x"27",   x"BE",   x"C9", 
  x"71",   x"06",   x"9F",   x"E8",   x"6E",   x"19",   x"80",   x"F7", 
  x"CB",   x"BC",   x"25",   x"52",   x"D4",   x"A3",   x"3A",   x"4D", 
  x"F5",   x"82",   x"1B",   x"6C",   x"EA",   x"9D",   x"04",   x"73", 
  x"B7",   x"C0",   x"59",   x"2E",   x"A8",   x"DF",   x"46",   x"31", 
  x"89",   x"FE",   x"67",   x"10",   x"96",   x"E1",   x"78",   x"0F", 
  x"66",   x"11",   x"88",   x"FF",   x"79",   x"0E",   x"97",   x"E0", 
  x"58",   x"2F",   x"B6",   x"C1",   x"47",   x"30",   x"A9",   x"DE", 
  x"1A",   x"6D",   x"F4",   x"83",   x"05",   x"72",   x"EB",   x"9C", 
  x"24",   x"53",   x"CA",   x"BD",   x"3B",   x"4C",   x"D5",   x"A2", 
  x"9E",   x"E9",   x"70",   x"07",   x"81",   x"F6",   x"6F",   x"18", 
  x"A0",   x"D7",   x"4E",   x"39",   x"BF",   x"C8",   x"51",   x"26", 
  x"E2",   x"95",   x"0C",   x"7B",   x"FD",   x"8A",   x"13",   x"64", 
  x"DC",   x"AB",   x"32",   x"45",   x"C3",   x"B4",   x"2D",   x"5A", 
  x"55",   x"22",   x"BB",   x"CC",   x"4A",   x"3D",   x"A4",   x"D3", 
  x"6B",   x"1C",   x"85",   x"F2",   x"74",   x"03",   x"9A",   x"ED", 
  x"29",   x"5E",   x"C7",   x"B0",   x"36",   x"41",   x"D8",   x"AF", 
  x"17",   x"60",   x"F9",   x"8E",   x"08",   x"7F",   x"E6",   x"91", 
  x"AD",   x"DA",   x"43",   x"34",   x"B2",   x"C5",   x"5C",   x"2B", 
  x"93",   x"E4",   x"7D",   x"0A",   x"8C",   x"FB",   x"62",   x"15", 
  x"D1",   x"A6",   x"3F",   x"48",   x"CE",   x"B9",   x"20",   x"57", 
  x"EF",   x"98",   x"01",   x"76",   x"F0",   x"87",   x"1E",   x"69", 
  x"00",   x"78",   x"F0",   x"88",   x"23",   x"5B",   x"D3",   x"AB", 
  x"46",   x"3E",   x"B6",   x"CE",   x"65",   x"1D",   x"95",   x"ED", 
  x"8C",   x"F4",   x"7C",   x"04",   x"AF",   x"D7",   x"5F",   x"27", 
  x"CA",   x"B2",   x"3A",   x"42",   x"E9",   x"91",   x"19",   x"61", 
  x"DB",   x"A3",   x"2B",   x"53",   x"F8",   x"80",   x"08",   x"70", 
  x"9D",   x"E5",   x"6D",   x"15",   x"BE",   x"C6",   x"4E",   x"36", 
  x"57",   x"2F",   x"A7",   x"DF",   x"74",   x"0C",   x"84",   x"FC", 
  x"11",   x"69",   x"E1",   x"99",   x"32",   x"4A",   x"C2",   x"BA", 
  x"75",   x"0D",   x"85",   x"FD",   x"56",   x"2E",   x"A6",   x"DE", 
  x"33",   x"4B",   x"C3",   x"BB",   x"10",   x"68",   x"E0",   x"98", 
  x"F9",   x"81",   x"09",   x"71",   x"DA",   x"A2",   x"2A",   x"52", 
  x"BF",   x"C7",   x"4F",   x"37",   x"9C",   x"E4",   x"6C",   x"14", 
  x"AE",   x"D6",   x"5E",   x"26",   x"8D",   x"F5",   x"7D",   x"05", 
  x"E8",   x"90",   x"18",   x"60",   x"CB",   x"B3",   x"3B",   x"43", 
  x"22",   x"5A",   x"D2",   x"AA",   x"01",   x"79",   x"F1",   x"89", 
  x"64",   x"1C",   x"94",   x"EC",   x"47",   x"3F",   x"B7",   x"CF", 
  x"EA",   x"92",   x"1A",   x"62",   x"C9",   x"B1",   x"39",   x"41", 
  x"AC",   x"D4",   x"5C",   x"24",   x"8F",   x"F7",   x"7F",   x"07", 
  x"66",   x"1E",   x"96",   x"EE",   x"45",   x"3D",   x"B5",   x"CD", 
  x"20",   x"58",   x"D0",   x"A8",   x"03",   x"7B",   x"F3",   x"8B", 
  x"31",   x"49",   x"C1",   x"B9",   x"12",   x"6A",   x"E2",   x"9A", 
  x"77",   x"0F",   x"87",   x"FF",   x"54",   x"2C",   x"A4",   x"DC", 
  x"BD",   x"C5",   x"4D",   x"35",   x"9E",   x"E6",   x"6E",   x"16", 
  x"FB",   x"83",   x"0B",   x"73",   x"D8",   x"A0",   x"28",   x"50", 
  x"9F",   x"E7",   x"6F",   x"17",   x"BC",   x"C4",   x"4C",   x"34", 
  x"D9",   x"A1",   x"29",   x"51",   x"FA",   x"82",   x"0A",   x"72", 
  x"13",   x"6B",   x"E3",   x"9B",   x"30",   x"48",   x"C0",   x"B8", 
  x"55",   x"2D",   x"A5",   x"DD",   x"76",   x"0E",   x"86",   x"FE", 
  x"44",   x"3C",   x"B4",   x"CC",   x"67",   x"1F",   x"97",   x"EF", 
  x"02",   x"7A",   x"F2",   x"8A",   x"21",   x"59",   x"D1",   x"A9", 
  x"C8",   x"B0",   x"38",   x"40",   x"EB",   x"93",   x"1B",   x"63", 
  x"8E",   x"F6",   x"7E",   x"06",   x"AD",   x"D5",   x"5D",   x"25", 
  x"00",   x"79",   x"F2",   x"8B",   x"27",   x"5E",   x"D5",   x"AC", 
  x"4E",   x"37",   x"BC",   x"C5",   x"69",   x"10",   x"9B",   x"E2", 
  x"9C",   x"E5",   x"6E",   x"17",   x"BB",   x"C2",   x"49",   x"30", 
  x"D2",   x"AB",   x"20",   x"59",   x"F5",   x"8C",   x"07",   x"7E", 
  x"FB",   x"82",   x"09",   x"70",   x"DC",   x"A5",   x"2E",   x"57", 
  x"B5",   x"CC",   x"47",   x"3E",   x"92",   x"EB",   x"60",   x"19", 
  x"67",   x"1E",   x"95",   x"EC",   x"40",   x"39",   x"B2",   x"CB", 
  x"29",   x"50",   x"DB",   x"A2",   x"0E",   x"77",   x"FC",   x"85", 
  x"35",   x"4C",   x"C7",   x"BE",   x"12",   x"6B",   x"E0",   x"99", 
  x"7B",   x"02",   x"89",   x"F0",   x"5C",   x"25",   x"AE",   x"D7", 
  x"A9",   x"D0",   x"5B",   x"22",   x"8E",   x"F7",   x"7C",   x"05", 
  x"E7",   x"9E",   x"15",   x"6C",   x"C0",   x"B9",   x"32",   x"4B", 
  x"CE",   x"B7",   x"3C",   x"45",   x"E9",   x"90",   x"1B",   x"62", 
  x"80",   x"F9",   x"72",   x"0B",   x"A7",   x"DE",   x"55",   x"2C", 
  x"52",   x"2B",   x"A0",   x"D9",   x"75",   x"0C",   x"87",   x"FE", 
  x"1C",   x"65",   x"EE",   x"97",   x"3B",   x"42",   x"C9",   x"B0", 
  x"6A",   x"13",   x"98",   x"E1",   x"4D",   x"34",   x"BF",   x"C6", 
  x"24",   x"5D",   x"D6",   x"AF",   x"03",   x"7A",   x"F1",   x"88", 
  x"F6",   x"8F",   x"04",   x"7D",   x"D1",   x"A8",   x"23",   x"5A", 
  x"B8",   x"C1",   x"4A",   x"33",   x"9F",   x"E6",   x"6D",   x"14", 
  x"91",   x"E8",   x"63",   x"1A",   x"B6",   x"CF",   x"44",   x"3D", 
  x"DF",   x"A6",   x"2D",   x"54",   x"F8",   x"81",   x"0A",   x"73", 
  x"0D",   x"74",   x"FF",   x"86",   x"2A",   x"53",   x"D8",   x"A1", 
  x"43",   x"3A",   x"B1",   x"C8",   x"64",   x"1D",   x"96",   x"EF", 
  x"5F",   x"26",   x"AD",   x"D4",   x"78",   x"01",   x"8A",   x"F3", 
  x"11",   x"68",   x"E3",   x"9A",   x"36",   x"4F",   x"C4",   x"BD", 
  x"C3",   x"BA",   x"31",   x"48",   x"E4",   x"9D",   x"16",   x"6F", 
  x"8D",   x"F4",   x"7F",   x"06",   x"AA",   x"D3",   x"58",   x"21", 
  x"A4",   x"DD",   x"56",   x"2F",   x"83",   x"FA",   x"71",   x"08", 
  x"EA",   x"93",   x"18",   x"61",   x"CD",   x"B4",   x"3F",   x"46", 
  x"38",   x"41",   x"CA",   x"B3",   x"1F",   x"66",   x"ED",   x"94", 
  x"76",   x"0F",   x"84",   x"FD",   x"51",   x"28",   x"A3",   x"DA", 
  x"00",   x"7A",   x"F4",   x"8E",   x"2B",   x"51",   x"DF",   x"A5", 
  x"56",   x"2C",   x"A2",   x"D8",   x"7D",   x"07",   x"89",   x"F3", 
  x"AC",   x"D6",   x"58",   x"22",   x"87",   x"FD",   x"73",   x"09", 
  x"FA",   x"80",   x"0E",   x"74",   x"D1",   x"AB",   x"25",   x"5F", 
  x"9B",   x"E1",   x"6F",   x"15",   x"B0",   x"CA",   x"44",   x"3E", 
  x"CD",   x"B7",   x"39",   x"43",   x"E6",   x"9C",   x"12",   x"68", 
  x"37",   x"4D",   x"C3",   x"B9",   x"1C",   x"66",   x"E8",   x"92", 
  x"61",   x"1B",   x"95",   x"EF",   x"4A",   x"30",   x"BE",   x"C4", 
  x"F5",   x"8F",   x"01",   x"7B",   x"DE",   x"A4",   x"2A",   x"50", 
  x"A3",   x"D9",   x"57",   x"2D",   x"88",   x"F2",   x"7C",   x"06", 
  x"59",   x"23",   x"AD",   x"D7",   x"72",   x"08",   x"86",   x"FC", 
  x"0F",   x"75",   x"FB",   x"81",   x"24",   x"5E",   x"D0",   x"AA", 
  x"6E",   x"14",   x"9A",   x"E0",   x"45",   x"3F",   x"B1",   x"CB", 
  x"38",   x"42",   x"CC",   x"B6",   x"13",   x"69",   x"E7",   x"9D", 
  x"C2",   x"B8",   x"36",   x"4C",   x"E9",   x"93",   x"1D",   x"67", 
  x"94",   x"EE",   x"60",   x"1A",   x"BF",   x"C5",   x"4B",   x"31", 
  x"29",   x"53",   x"DD",   x"A7",   x"02",   x"78",   x"F6",   x"8C", 
  x"7F",   x"05",   x"8B",   x"F1",   x"54",   x"2E",   x"A0",   x"DA", 
  x"85",   x"FF",   x"71",   x"0B",   x"AE",   x"D4",   x"5A",   x"20", 
  x"D3",   x"A9",   x"27",   x"5D",   x"F8",   x"82",   x"0C",   x"76", 
  x"B2",   x"C8",   x"46",   x"3C",   x"99",   x"E3",   x"6D",   x"17", 
  x"E4",   x"9E",   x"10",   x"6A",   x"CF",   x"B5",   x"3B",   x"41", 
  x"1E",   x"64",   x"EA",   x"90",   x"35",   x"4F",   x"C1",   x"BB", 
  x"48",   x"32",   x"BC",   x"C6",   x"63",   x"19",   x"97",   x"ED", 
  x"DC",   x"A6",   x"28",   x"52",   x"F7",   x"8D",   x"03",   x"79", 
  x"8A",   x"F0",   x"7E",   x"04",   x"A1",   x"DB",   x"55",   x"2F", 
  x"70",   x"0A",   x"84",   x"FE",   x"5B",   x"21",   x"AF",   x"D5", 
  x"26",   x"5C",   x"D2",   x"A8",   x"0D",   x"77",   x"F9",   x"83", 
  x"47",   x"3D",   x"B3",   x"C9",   x"6C",   x"16",   x"98",   x"E2", 
  x"11",   x"6B",   x"E5",   x"9F",   x"3A",   x"40",   x"CE",   x"B4", 
  x"EB",   x"91",   x"1F",   x"65",   x"C0",   x"BA",   x"34",   x"4E", 
  x"BD",   x"C7",   x"49",   x"33",   x"96",   x"EC",   x"62",   x"18", 
  x"00",   x"7B",   x"F6",   x"8D",   x"2F",   x"54",   x"D9",   x"A2", 
  x"5E",   x"25",   x"A8",   x"D3",   x"71",   x"0A",   x"87",   x"FC", 
  x"BC",   x"C7",   x"4A",   x"31",   x"93",   x"E8",   x"65",   x"1E", 
  x"E2",   x"99",   x"14",   x"6F",   x"CD",   x"B6",   x"3B",   x"40", 
  x"BB",   x"C0",   x"4D",   x"36",   x"94",   x"EF",   x"62",   x"19", 
  x"E5",   x"9E",   x"13",   x"68",   x"CA",   x"B1",   x"3C",   x"47", 
  x"07",   x"7C",   x"F1",   x"8A",   x"28",   x"53",   x"DE",   x"A5", 
  x"59",   x"22",   x"AF",   x"D4",   x"76",   x"0D",   x"80",   x"FB", 
  x"B5",   x"CE",   x"43",   x"38",   x"9A",   x"E1",   x"6C",   x"17", 
  x"EB",   x"90",   x"1D",   x"66",   x"C4",   x"BF",   x"32",   x"49", 
  x"09",   x"72",   x"FF",   x"84",   x"26",   x"5D",   x"D0",   x"AB", 
  x"57",   x"2C",   x"A1",   x"DA",   x"78",   x"03",   x"8E",   x"F5", 
  x"0E",   x"75",   x"F8",   x"83",   x"21",   x"5A",   x"D7",   x"AC", 
  x"50",   x"2B",   x"A6",   x"DD",   x"7F",   x"04",   x"89",   x"F2", 
  x"B2",   x"C9",   x"44",   x"3F",   x"9D",   x"E6",   x"6B",   x"10", 
  x"EC",   x"97",   x"1A",   x"61",   x"C3",   x"B8",   x"35",   x"4E", 
  x"A9",   x"D2",   x"5F",   x"24",   x"86",   x"FD",   x"70",   x"0B", 
  x"F7",   x"8C",   x"01",   x"7A",   x"D8",   x"A3",   x"2E",   x"55", 
  x"15",   x"6E",   x"E3",   x"98",   x"3A",   x"41",   x"CC",   x"B7", 
  x"4B",   x"30",   x"BD",   x"C6",   x"64",   x"1F",   x"92",   x"E9", 
  x"12",   x"69",   x"E4",   x"9F",   x"3D",   x"46",   x"CB",   x"B0", 
  x"4C",   x"37",   x"BA",   x"C1",   x"63",   x"18",   x"95",   x"EE", 
  x"AE",   x"D5",   x"58",   x"23",   x"81",   x"FA",   x"77",   x"0C", 
  x"F0",   x"8B",   x"06",   x"7D",   x"DF",   x"A4",   x"29",   x"52", 
  x"1C",   x"67",   x"EA",   x"91",   x"33",   x"48",   x"C5",   x"BE", 
  x"42",   x"39",   x"B4",   x"CF",   x"6D",   x"16",   x"9B",   x"E0", 
  x"A0",   x"DB",   x"56",   x"2D",   x"8F",   x"F4",   x"79",   x"02", 
  x"FE",   x"85",   x"08",   x"73",   x"D1",   x"AA",   x"27",   x"5C", 
  x"A7",   x"DC",   x"51",   x"2A",   x"88",   x"F3",   x"7E",   x"05", 
  x"F9",   x"82",   x"0F",   x"74",   x"D6",   x"AD",   x"20",   x"5B", 
  x"1B",   x"60",   x"ED",   x"96",   x"34",   x"4F",   x"C2",   x"B9", 
  x"45",   x"3E",   x"B3",   x"C8",   x"6A",   x"11",   x"9C",   x"E7", 
  x"00",   x"7C",   x"F8",   x"84",   x"33",   x"4F",   x"CB",   x"B7", 
  x"66",   x"1A",   x"9E",   x"E2",   x"55",   x"29",   x"AD",   x"D1", 
  x"CC",   x"B0",   x"34",   x"48",   x"FF",   x"83",   x"07",   x"7B", 
  x"AA",   x"D6",   x"52",   x"2E",   x"99",   x"E5",   x"61",   x"1D", 
  x"5B",   x"27",   x"A3",   x"DF",   x"68",   x"14",   x"90",   x"EC", 
  x"3D",   x"41",   x"C5",   x"B9",   x"0E",   x"72",   x"F6",   x"8A", 
  x"97",   x"EB",   x"6F",   x"13",   x"A4",   x"D8",   x"5C",   x"20", 
  x"F1",   x"8D",   x"09",   x"75",   x"C2",   x"BE",   x"3A",   x"46", 
  x"B6",   x"CA",   x"4E",   x"32",   x"85",   x"F9",   x"7D",   x"01", 
  x"D0",   x"AC",   x"28",   x"54",   x"E3",   x"9F",   x"1B",   x"67", 
  x"7A",   x"06",   x"82",   x"FE",   x"49",   x"35",   x"B1",   x"CD", 
  x"1C",   x"60",   x"E4",   x"98",   x"2F",   x"53",   x"D7",   x"AB", 
  x"ED",   x"91",   x"15",   x"69",   x"DE",   x"A2",   x"26",   x"5A", 
  x"8B",   x"F7",   x"73",   x"0F",   x"B8",   x"C4",   x"40",   x"3C", 
  x"21",   x"5D",   x"D9",   x"A5",   x"12",   x"6E",   x"EA",   x"96", 
  x"47",   x"3B",   x"BF",   x"C3",   x"74",   x"08",   x"8C",   x"F0", 
  x"AF",   x"D3",   x"57",   x"2B",   x"9C",   x"E0",   x"64",   x"18", 
  x"C9",   x"B5",   x"31",   x"4D",   x"FA",   x"86",   x"02",   x"7E", 
  x"63",   x"1F",   x"9B",   x"E7",   x"50",   x"2C",   x"A8",   x"D4", 
  x"05",   x"79",   x"FD",   x"81",   x"36",   x"4A",   x"CE",   x"B2", 
  x"F4",   x"88",   x"0C",   x"70",   x"C7",   x"BB",   x"3F",   x"43", 
  x"92",   x"EE",   x"6A",   x"16",   x"A1",   x"DD",   x"59",   x"25", 
  x"38",   x"44",   x"C0",   x"BC",   x"0B",   x"77",   x"F3",   x"8F", 
  x"5E",   x"22",   x"A6",   x"DA",   x"6D",   x"11",   x"95",   x"E9", 
  x"19",   x"65",   x"E1",   x"9D",   x"2A",   x"56",   x"D2",   x"AE", 
  x"7F",   x"03",   x"87",   x"FB",   x"4C",   x"30",   x"B4",   x"C8", 
  x"D5",   x"A9",   x"2D",   x"51",   x"E6",   x"9A",   x"1E",   x"62", 
  x"B3",   x"CF",   x"4B",   x"37",   x"80",   x"FC",   x"78",   x"04", 
  x"42",   x"3E",   x"BA",   x"C6",   x"71",   x"0D",   x"89",   x"F5", 
  x"24",   x"58",   x"DC",   x"A0",   x"17",   x"6B",   x"EF",   x"93", 
  x"8E",   x"F2",   x"76",   x"0A",   x"BD",   x"C1",   x"45",   x"39", 
  x"E8",   x"94",   x"10",   x"6C",   x"DB",   x"A7",   x"23",   x"5F", 
  x"00",   x"7D",   x"FA",   x"87",   x"37",   x"4A",   x"CD",   x"B0", 
  x"6E",   x"13",   x"94",   x"E9",   x"59",   x"24",   x"A3",   x"DE", 
  x"DC",   x"A1",   x"26",   x"5B",   x"EB",   x"96",   x"11",   x"6C", 
  x"B2",   x"CF",   x"48",   x"35",   x"85",   x"F8",   x"7F",   x"02", 
  x"7B",   x"06",   x"81",   x"FC",   x"4C",   x"31",   x"B6",   x"CB", 
  x"15",   x"68",   x"EF",   x"92",   x"22",   x"5F",   x"D8",   x"A5", 
  x"A7",   x"DA",   x"5D",   x"20",   x"90",   x"ED",   x"6A",   x"17", 
  x"C9",   x"B4",   x"33",   x"4E",   x"FE",   x"83",   x"04",   x"79", 
  x"F6",   x"8B",   x"0C",   x"71",   x"C1",   x"BC",   x"3B",   x"46", 
  x"98",   x"E5",   x"62",   x"1F",   x"AF",   x"D2",   x"55",   x"28", 
  x"2A",   x"57",   x"D0",   x"AD",   x"1D",   x"60",   x"E7",   x"9A", 
  x"44",   x"39",   x"BE",   x"C3",   x"73",   x"0E",   x"89",   x"F4", 
  x"8D",   x"F0",   x"77",   x"0A",   x"BA",   x"C7",   x"40",   x"3D", 
  x"E3",   x"9E",   x"19",   x"64",   x"D4",   x"A9",   x"2E",   x"53", 
  x"51",   x"2C",   x"AB",   x"D6",   x"66",   x"1B",   x"9C",   x"E1", 
  x"3F",   x"42",   x"C5",   x"B8",   x"08",   x"75",   x"F2",   x"8F", 
  x"2F",   x"52",   x"D5",   x"A8",   x"18",   x"65",   x"E2",   x"9F", 
  x"41",   x"3C",   x"BB",   x"C6",   x"76",   x"0B",   x"8C",   x"F1", 
  x"F3",   x"8E",   x"09",   x"74",   x"C4",   x"B9",   x"3E",   x"43", 
  x"9D",   x"E0",   x"67",   x"1A",   x"AA",   x"D7",   x"50",   x"2D", 
  x"54",   x"29",   x"AE",   x"D3",   x"63",   x"1E",   x"99",   x"E4", 
  x"3A",   x"47",   x"C0",   x"BD",   x"0D",   x"70",   x"F7",   x"8A", 
  x"88",   x"F5",   x"72",   x"0F",   x"BF",   x"C2",   x"45",   x"38", 
  x"E6",   x"9B",   x"1C",   x"61",   x"D1",   x"AC",   x"2B",   x"56", 
  x"D9",   x"A4",   x"23",   x"5E",   x"EE",   x"93",   x"14",   x"69", 
  x"B7",   x"CA",   x"4D",   x"30",   x"80",   x"FD",   x"7A",   x"07", 
  x"05",   x"78",   x"FF",   x"82",   x"32",   x"4F",   x"C8",   x"B5", 
  x"6B",   x"16",   x"91",   x"EC",   x"5C",   x"21",   x"A6",   x"DB", 
  x"A2",   x"DF",   x"58",   x"25",   x"95",   x"E8",   x"6F",   x"12", 
  x"CC",   x"B1",   x"36",   x"4B",   x"FB",   x"86",   x"01",   x"7C", 
  x"7E",   x"03",   x"84",   x"F9",   x"49",   x"34",   x"B3",   x"CE", 
  x"10",   x"6D",   x"EA",   x"97",   x"27",   x"5A",   x"DD",   x"A0", 
  x"00",   x"7E",   x"FC",   x"82",   x"3B",   x"45",   x"C7",   x"B9", 
  x"76",   x"08",   x"8A",   x"F4",   x"4D",   x"33",   x"B1",   x"CF", 
  x"EC",   x"92",   x"10",   x"6E",   x"D7",   x"A9",   x"2B",   x"55", 
  x"9A",   x"E4",   x"66",   x"18",   x"A1",   x"DF",   x"5D",   x"23", 
  x"1B",   x"65",   x"E7",   x"99",   x"20",   x"5E",   x"DC",   x"A2", 
  x"6D",   x"13",   x"91",   x"EF",   x"56",   x"28",   x"AA",   x"D4", 
  x"F7",   x"89",   x"0B",   x"75",   x"CC",   x"B2",   x"30",   x"4E", 
  x"81",   x"FF",   x"7D",   x"03",   x"BA",   x"C4",   x"46",   x"38", 
  x"36",   x"48",   x"CA",   x"B4",   x"0D",   x"73",   x"F1",   x"8F", 
  x"40",   x"3E",   x"BC",   x"C2",   x"7B",   x"05",   x"87",   x"F9", 
  x"DA",   x"A4",   x"26",   x"58",   x"E1",   x"9F",   x"1D",   x"63", 
  x"AC",   x"D2",   x"50",   x"2E",   x"97",   x"E9",   x"6B",   x"15", 
  x"2D",   x"53",   x"D1",   x"AF",   x"16",   x"68",   x"EA",   x"94", 
  x"5B",   x"25",   x"A7",   x"D9",   x"60",   x"1E",   x"9C",   x"E2", 
  x"C1",   x"BF",   x"3D",   x"43",   x"FA",   x"84",   x"06",   x"78", 
  x"B7",   x"C9",   x"4B",   x"35",   x"8C",   x"F2",   x"70",   x"0E", 
  x"6C",   x"12",   x"90",   x"EE",   x"57",   x"29",   x"AB",   x"D5", 
  x"1A",   x"64",   x"E6",   x"98",   x"21",   x"5F",   x"DD",   x"A3", 
  x"80",   x"FE",   x"7C",   x"02",   x"BB",   x"C5",   x"47",   x"39", 
  x"F6",   x"88",   x"0A",   x"74",   x"CD",   x"B3",   x"31",   x"4F", 
  x"77",   x"09",   x"8B",   x"F5",   x"4C",   x"32",   x"B0",   x"CE", 
  x"01",   x"7F",   x"FD",   x"83",   x"3A",   x"44",   x"C6",   x"B8", 
  x"9B",   x"E5",   x"67",   x"19",   x"A0",   x"DE",   x"5C",   x"22", 
  x"ED",   x"93",   x"11",   x"6F",   x"D6",   x"A8",   x"2A",   x"54", 
  x"5A",   x"24",   x"A6",   x"D8",   x"61",   x"1F",   x"9D",   x"E3", 
  x"2C",   x"52",   x"D0",   x"AE",   x"17",   x"69",   x"EB",   x"95", 
  x"B6",   x"C8",   x"4A",   x"34",   x"8D",   x"F3",   x"71",   x"0F", 
  x"C0",   x"BE",   x"3C",   x"42",   x"FB",   x"85",   x"07",   x"79", 
  x"41",   x"3F",   x"BD",   x"C3",   x"7A",   x"04",   x"86",   x"F8", 
  x"37",   x"49",   x"CB",   x"B5",   x"0C",   x"72",   x"F0",   x"8E", 
  x"AD",   x"D3",   x"51",   x"2F",   x"96",   x"E8",   x"6A",   x"14", 
  x"DB",   x"A5",   x"27",   x"59",   x"E0",   x"9E",   x"1C",   x"62", 
  x"00",   x"7F",   x"FE",   x"81",   x"3F",   x"40",   x"C1",   x"BE", 
  x"7E",   x"01",   x"80",   x"FF",   x"41",   x"3E",   x"BF",   x"C0", 
  x"FC",   x"83",   x"02",   x"7D",   x"C3",   x"BC",   x"3D",   x"42", 
  x"82",   x"FD",   x"7C",   x"03",   x"BD",   x"C2",   x"43",   x"3C", 
  x"3B",   x"44",   x"C5",   x"BA",   x"04",   x"7B",   x"FA",   x"85", 
  x"45",   x"3A",   x"BB",   x"C4",   x"7A",   x"05",   x"84",   x"FB", 
  x"C7",   x"B8",   x"39",   x"46",   x"F8",   x"87",   x"06",   x"79", 
  x"B9",   x"C6",   x"47",   x"38",   x"86",   x"F9",   x"78",   x"07", 
  x"76",   x"09",   x"88",   x"F7",   x"49",   x"36",   x"B7",   x"C8", 
  x"08",   x"77",   x"F6",   x"89",   x"37",   x"48",   x"C9",   x"B6", 
  x"8A",   x"F5",   x"74",   x"0B",   x"B5",   x"CA",   x"4B",   x"34", 
  x"F4",   x"8B",   x"0A",   x"75",   x"CB",   x"B4",   x"35",   x"4A", 
  x"4D",   x"32",   x"B3",   x"CC",   x"72",   x"0D",   x"8C",   x"F3", 
  x"33",   x"4C",   x"CD",   x"B2",   x"0C",   x"73",   x"F2",   x"8D", 
  x"B1",   x"CE",   x"4F",   x"30",   x"8E",   x"F1",   x"70",   x"0F", 
  x"CF",   x"B0",   x"31",   x"4E",   x"F0",   x"8F",   x"0E",   x"71", 
  x"EC",   x"93",   x"12",   x"6D",   x"D3",   x"AC",   x"2D",   x"52", 
  x"92",   x"ED",   x"6C",   x"13",   x"AD",   x"D2",   x"53",   x"2C", 
  x"10",   x"6F",   x"EE",   x"91",   x"2F",   x"50",   x"D1",   x"AE", 
  x"6E",   x"11",   x"90",   x"EF",   x"51",   x"2E",   x"AF",   x"D0", 
  x"D7",   x"A8",   x"29",   x"56",   x"E8",   x"97",   x"16",   x"69", 
  x"A9",   x"D6",   x"57",   x"28",   x"96",   x"E9",   x"68",   x"17", 
  x"2B",   x"54",   x"D5",   x"AA",   x"14",   x"6B",   x"EA",   x"95", 
  x"55",   x"2A",   x"AB",   x"D4",   x"6A",   x"15",   x"94",   x"EB", 
  x"9A",   x"E5",   x"64",   x"1B",   x"A5",   x"DA",   x"5B",   x"24", 
  x"E4",   x"9B",   x"1A",   x"65",   x"DB",   x"A4",   x"25",   x"5A", 
  x"66",   x"19",   x"98",   x"E7",   x"59",   x"26",   x"A7",   x"D8", 
  x"18",   x"67",   x"E6",   x"99",   x"27",   x"58",   x"D9",   x"A6", 
  x"A1",   x"DE",   x"5F",   x"20",   x"9E",   x"E1",   x"60",   x"1F", 
  x"DF",   x"A0",   x"21",   x"5E",   x"E0",   x"9F",   x"1E",   x"61", 
  x"5D",   x"22",   x"A3",   x"DC",   x"62",   x"1D",   x"9C",   x"E3", 
  x"23",   x"5C",   x"DD",   x"A2",   x"1C",   x"63",   x"E2",   x"9D", 
  x"00",   x"80",   x"C3",   x"43",   x"45",   x"C5",   x"86",   x"06", 
  x"8A",   x"0A",   x"49",   x"C9",   x"CF",   x"4F",   x"0C",   x"8C", 
  x"D7",   x"57",   x"14",   x"94",   x"92",   x"12",   x"51",   x"D1", 
  x"5D",   x"DD",   x"9E",   x"1E",   x"18",   x"98",   x"DB",   x"5B", 
  x"6D",   x"ED",   x"AE",   x"2E",   x"28",   x"A8",   x"EB",   x"6B", 
  x"E7",   x"67",   x"24",   x"A4",   x"A2",   x"22",   x"61",   x"E1", 
  x"BA",   x"3A",   x"79",   x"F9",   x"FF",   x"7F",   x"3C",   x"BC", 
  x"30",   x"B0",   x"F3",   x"73",   x"75",   x"F5",   x"B6",   x"36", 
  x"DA",   x"5A",   x"19",   x"99",   x"9F",   x"1F",   x"5C",   x"DC", 
  x"50",   x"D0",   x"93",   x"13",   x"15",   x"95",   x"D6",   x"56", 
  x"0D",   x"8D",   x"CE",   x"4E",   x"48",   x"C8",   x"8B",   x"0B", 
  x"87",   x"07",   x"44",   x"C4",   x"C2",   x"42",   x"01",   x"81", 
  x"B7",   x"37",   x"74",   x"F4",   x"F2",   x"72",   x"31",   x"B1", 
  x"3D",   x"BD",   x"FE",   x"7E",   x"78",   x"F8",   x"BB",   x"3B", 
  x"60",   x"E0",   x"A3",   x"23",   x"25",   x"A5",   x"E6",   x"66", 
  x"EA",   x"6A",   x"29",   x"A9",   x"AF",   x"2F",   x"6C",   x"EC", 
  x"77",   x"F7",   x"B4",   x"34",   x"32",   x"B2",   x"F1",   x"71", 
  x"FD",   x"7D",   x"3E",   x"BE",   x"B8",   x"38",   x"7B",   x"FB", 
  x"A0",   x"20",   x"63",   x"E3",   x"E5",   x"65",   x"26",   x"A6", 
  x"2A",   x"AA",   x"E9",   x"69",   x"6F",   x"EF",   x"AC",   x"2C", 
  x"1A",   x"9A",   x"D9",   x"59",   x"5F",   x"DF",   x"9C",   x"1C", 
  x"90",   x"10",   x"53",   x"D3",   x"D5",   x"55",   x"16",   x"96", 
  x"CD",   x"4D",   x"0E",   x"8E",   x"88",   x"08",   x"4B",   x"CB", 
  x"47",   x"C7",   x"84",   x"04",   x"02",   x"82",   x"C1",   x"41", 
  x"AD",   x"2D",   x"6E",   x"EE",   x"E8",   x"68",   x"2B",   x"AB", 
  x"27",   x"A7",   x"E4",   x"64",   x"62",   x"E2",   x"A1",   x"21", 
  x"7A",   x"FA",   x"B9",   x"39",   x"3F",   x"BF",   x"FC",   x"7C", 
  x"F0",   x"70",   x"33",   x"B3",   x"B5",   x"35",   x"76",   x"F6", 
  x"C0",   x"40",   x"03",   x"83",   x"85",   x"05",   x"46",   x"C6", 
  x"4A",   x"CA",   x"89",   x"09",   x"0F",   x"8F",   x"CC",   x"4C", 
  x"17",   x"97",   x"D4",   x"54",   x"52",   x"D2",   x"91",   x"11", 
  x"9D",   x"1D",   x"5E",   x"DE",   x"D8",   x"58",   x"1B",   x"9B", 
  x"00",   x"81",   x"C1",   x"40",   x"41",   x"C0",   x"80",   x"01", 
  x"82",   x"03",   x"43",   x"C2",   x"C3",   x"42",   x"02",   x"83", 
  x"C7",   x"46",   x"06",   x"87",   x"86",   x"07",   x"47",   x"C6", 
  x"45",   x"C4",   x"84",   x"05",   x"04",   x"85",   x"C5",   x"44", 
  x"4D",   x"CC",   x"8C",   x"0D",   x"0C",   x"8D",   x"CD",   x"4C", 
  x"CF",   x"4E",   x"0E",   x"8F",   x"8E",   x"0F",   x"4F",   x"CE", 
  x"8A",   x"0B",   x"4B",   x"CA",   x"CB",   x"4A",   x"0A",   x"8B", 
  x"08",   x"89",   x"C9",   x"48",   x"49",   x"C8",   x"88",   x"09", 
  x"9A",   x"1B",   x"5B",   x"DA",   x"DB",   x"5A",   x"1A",   x"9B", 
  x"18",   x"99",   x"D9",   x"58",   x"59",   x"D8",   x"98",   x"19", 
  x"5D",   x"DC",   x"9C",   x"1D",   x"1C",   x"9D",   x"DD",   x"5C", 
  x"DF",   x"5E",   x"1E",   x"9F",   x"9E",   x"1F",   x"5F",   x"DE", 
  x"D7",   x"56",   x"16",   x"97",   x"96",   x"17",   x"57",   x"D6", 
  x"55",   x"D4",   x"94",   x"15",   x"14",   x"95",   x"D5",   x"54", 
  x"10",   x"91",   x"D1",   x"50",   x"51",   x"D0",   x"90",   x"11", 
  x"92",   x"13",   x"53",   x"D2",   x"D3",   x"52",   x"12",   x"93", 
  x"F7",   x"76",   x"36",   x"B7",   x"B6",   x"37",   x"77",   x"F6", 
  x"75",   x"F4",   x"B4",   x"35",   x"34",   x"B5",   x"F5",   x"74", 
  x"30",   x"B1",   x"F1",   x"70",   x"71",   x"F0",   x"B0",   x"31", 
  x"B2",   x"33",   x"73",   x"F2",   x"F3",   x"72",   x"32",   x"B3", 
  x"BA",   x"3B",   x"7B",   x"FA",   x"FB",   x"7A",   x"3A",   x"BB", 
  x"38",   x"B9",   x"F9",   x"78",   x"79",   x"F8",   x"B8",   x"39", 
  x"7D",   x"FC",   x"BC",   x"3D",   x"3C",   x"BD",   x"FD",   x"7C", 
  x"FF",   x"7E",   x"3E",   x"BF",   x"BE",   x"3F",   x"7F",   x"FE", 
  x"6D",   x"EC",   x"AC",   x"2D",   x"2C",   x"AD",   x"ED",   x"6C", 
  x"EF",   x"6E",   x"2E",   x"AF",   x"AE",   x"2F",   x"6F",   x"EE", 
  x"AA",   x"2B",   x"6B",   x"EA",   x"EB",   x"6A",   x"2A",   x"AB", 
  x"28",   x"A9",   x"E9",   x"68",   x"69",   x"E8",   x"A8",   x"29", 
  x"20",   x"A1",   x"E1",   x"60",   x"61",   x"E0",   x"A0",   x"21", 
  x"A2",   x"23",   x"63",   x"E2",   x"E3",   x"62",   x"22",   x"A3", 
  x"E7",   x"66",   x"26",   x"A7",   x"A6",   x"27",   x"67",   x"E6", 
  x"65",   x"E4",   x"A4",   x"25",   x"24",   x"A5",   x"E5",   x"64", 
  x"00",   x"82",   x"C7",   x"45",   x"4D",   x"CF",   x"8A",   x"08", 
  x"9A",   x"18",   x"5D",   x"DF",   x"D7",   x"55",   x"10",   x"92", 
  x"F7",   x"75",   x"30",   x"B2",   x"BA",   x"38",   x"7D",   x"FF", 
  x"6D",   x"EF",   x"AA",   x"28",   x"20",   x"A2",   x"E7",   x"65", 
  x"2D",   x"AF",   x"EA",   x"68",   x"60",   x"E2",   x"A7",   x"25", 
  x"B7",   x"35",   x"70",   x"F2",   x"FA",   x"78",   x"3D",   x"BF", 
  x"DA",   x"58",   x"1D",   x"9F",   x"97",   x"15",   x"50",   x"D2", 
  x"40",   x"C2",   x"87",   x"05",   x"0D",   x"8F",   x"CA",   x"48", 
  x"5A",   x"D8",   x"9D",   x"1F",   x"17",   x"95",   x"D0",   x"52", 
  x"C0",   x"42",   x"07",   x"85",   x"8D",   x"0F",   x"4A",   x"C8", 
  x"AD",   x"2F",   x"6A",   x"E8",   x"E0",   x"62",   x"27",   x"A5", 
  x"37",   x"B5",   x"F0",   x"72",   x"7A",   x"F8",   x"BD",   x"3F", 
  x"77",   x"F5",   x"B0",   x"32",   x"3A",   x"B8",   x"FD",   x"7F", 
  x"ED",   x"6F",   x"2A",   x"A8",   x"A0",   x"22",   x"67",   x"E5", 
  x"80",   x"02",   x"47",   x"C5",   x"CD",   x"4F",   x"0A",   x"88", 
  x"1A",   x"98",   x"DD",   x"5F",   x"57",   x"D5",   x"90",   x"12", 
  x"B4",   x"36",   x"73",   x"F1",   x"F9",   x"7B",   x"3E",   x"BC", 
  x"2E",   x"AC",   x"E9",   x"6B",   x"63",   x"E1",   x"A4",   x"26", 
  x"43",   x"C1",   x"84",   x"06",   x"0E",   x"8C",   x"C9",   x"4B", 
  x"D9",   x"5B",   x"1E",   x"9C",   x"94",   x"16",   x"53",   x"D1", 
  x"99",   x"1B",   x"5E",   x"DC",   x"D4",   x"56",   x"13",   x"91", 
  x"03",   x"81",   x"C4",   x"46",   x"4E",   x"CC",   x"89",   x"0B", 
  x"6E",   x"EC",   x"A9",   x"2B",   x"23",   x"A1",   x"E4",   x"66", 
  x"F4",   x"76",   x"33",   x"B1",   x"B9",   x"3B",   x"7E",   x"FC", 
  x"EE",   x"6C",   x"29",   x"AB",   x"A3",   x"21",   x"64",   x"E6", 
  x"74",   x"F6",   x"B3",   x"31",   x"39",   x"BB",   x"FE",   x"7C", 
  x"19",   x"9B",   x"DE",   x"5C",   x"54",   x"D6",   x"93",   x"11", 
  x"83",   x"01",   x"44",   x"C6",   x"CE",   x"4C",   x"09",   x"8B", 
  x"C3",   x"41",   x"04",   x"86",   x"8E",   x"0C",   x"49",   x"CB", 
  x"59",   x"DB",   x"9E",   x"1C",   x"14",   x"96",   x"D3",   x"51", 
  x"34",   x"B6",   x"F3",   x"71",   x"79",   x"FB",   x"BE",   x"3C", 
  x"AE",   x"2C",   x"69",   x"EB",   x"E3",   x"61",   x"24",   x"A6", 
  x"00",   x"83",   x"C5",   x"46",   x"49",   x"CA",   x"8C",   x"0F", 
  x"92",   x"11",   x"57",   x"D4",   x"DB",   x"58",   x"1E",   x"9D", 
  x"E7",   x"64",   x"22",   x"A1",   x"AE",   x"2D",   x"6B",   x"E8", 
  x"75",   x"F6",   x"B0",   x"33",   x"3C",   x"BF",   x"F9",   x"7A", 
  x"0D",   x"8E",   x"C8",   x"4B",   x"44",   x"C7",   x"81",   x"02", 
  x"9F",   x"1C",   x"5A",   x"D9",   x"D6",   x"55",   x"13",   x"90", 
  x"EA",   x"69",   x"2F",   x"AC",   x"A3",   x"20",   x"66",   x"E5", 
  x"78",   x"FB",   x"BD",   x"3E",   x"31",   x"B2",   x"F4",   x"77", 
  x"1A",   x"99",   x"DF",   x"5C",   x"53",   x"D0",   x"96",   x"15", 
  x"88",   x"0B",   x"4D",   x"CE",   x"C1",   x"42",   x"04",   x"87", 
  x"FD",   x"7E",   x"38",   x"BB",   x"B4",   x"37",   x"71",   x"F2", 
  x"6F",   x"EC",   x"AA",   x"29",   x"26",   x"A5",   x"E3",   x"60", 
  x"17",   x"94",   x"D2",   x"51",   x"5E",   x"DD",   x"9B",   x"18", 
  x"85",   x"06",   x"40",   x"C3",   x"CC",   x"4F",   x"09",   x"8A", 
  x"F0",   x"73",   x"35",   x"B6",   x"B9",   x"3A",   x"7C",   x"FF", 
  x"62",   x"E1",   x"A7",   x"24",   x"2B",   x"A8",   x"EE",   x"6D", 
  x"34",   x"B7",   x"F1",   x"72",   x"7D",   x"FE",   x"B8",   x"3B", 
  x"A6",   x"25",   x"63",   x"E0",   x"EF",   x"6C",   x"2A",   x"A9", 
  x"D3",   x"50",   x"16",   x"95",   x"9A",   x"19",   x"5F",   x"DC", 
  x"41",   x"C2",   x"84",   x"07",   x"08",   x"8B",   x"CD",   x"4E", 
  x"39",   x"BA",   x"FC",   x"7F",   x"70",   x"F3",   x"B5",   x"36", 
  x"AB",   x"28",   x"6E",   x"ED",   x"E2",   x"61",   x"27",   x"A4", 
  x"DE",   x"5D",   x"1B",   x"98",   x"97",   x"14",   x"52",   x"D1", 
  x"4C",   x"CF",   x"89",   x"0A",   x"05",   x"86",   x"C0",   x"43", 
  x"2E",   x"AD",   x"EB",   x"68",   x"67",   x"E4",   x"A2",   x"21", 
  x"BC",   x"3F",   x"79",   x"FA",   x"F5",   x"76",   x"30",   x"B3", 
  x"C9",   x"4A",   x"0C",   x"8F",   x"80",   x"03",   x"45",   x"C6", 
  x"5B",   x"D8",   x"9E",   x"1D",   x"12",   x"91",   x"D7",   x"54", 
  x"23",   x"A0",   x"E6",   x"65",   x"6A",   x"E9",   x"AF",   x"2C", 
  x"B1",   x"32",   x"74",   x"F7",   x"F8",   x"7B",   x"3D",   x"BE", 
  x"C4",   x"47",   x"01",   x"82",   x"8D",   x"0E",   x"48",   x"CB", 
  x"56",   x"D5",   x"93",   x"10",   x"1F",   x"9C",   x"DA",   x"59", 
  x"00",   x"84",   x"CB",   x"4F",   x"55",   x"D1",   x"9E",   x"1A", 
  x"AA",   x"2E",   x"61",   x"E5",   x"FF",   x"7B",   x"34",   x"B0", 
  x"97",   x"13",   x"5C",   x"D8",   x"C2",   x"46",   x"09",   x"8D", 
  x"3D",   x"B9",   x"F6",   x"72",   x"68",   x"EC",   x"A3",   x"27", 
  x"ED",   x"69",   x"26",   x"A2",   x"B8",   x"3C",   x"73",   x"F7", 
  x"47",   x"C3",   x"8C",   x"08",   x"12",   x"96",   x"D9",   x"5D", 
  x"7A",   x"FE",   x"B1",   x"35",   x"2F",   x"AB",   x"E4",   x"60", 
  x"D0",   x"54",   x"1B",   x"9F",   x"85",   x"01",   x"4E",   x"CA", 
  x"19",   x"9D",   x"D2",   x"56",   x"4C",   x"C8",   x"87",   x"03", 
  x"B3",   x"37",   x"78",   x"FC",   x"E6",   x"62",   x"2D",   x"A9", 
  x"8E",   x"0A",   x"45",   x"C1",   x"DB",   x"5F",   x"10",   x"94", 
  x"24",   x"A0",   x"EF",   x"6B",   x"71",   x"F5",   x"BA",   x"3E", 
  x"F4",   x"70",   x"3F",   x"BB",   x"A1",   x"25",   x"6A",   x"EE", 
  x"5E",   x"DA",   x"95",   x"11",   x"0B",   x"8F",   x"C0",   x"44", 
  x"63",   x"E7",   x"A8",   x"2C",   x"36",   x"B2",   x"FD",   x"79", 
  x"C9",   x"4D",   x"02",   x"86",   x"9C",   x"18",   x"57",   x"D3", 
  x"32",   x"B6",   x"F9",   x"7D",   x"67",   x"E3",   x"AC",   x"28", 
  x"98",   x"1C",   x"53",   x"D7",   x"CD",   x"49",   x"06",   x"82", 
  x"A5",   x"21",   x"6E",   x"EA",   x"F0",   x"74",   x"3B",   x"BF", 
  x"0F",   x"8B",   x"C4",   x"40",   x"5A",   x"DE",   x"91",   x"15", 
  x"DF",   x"5B",   x"14",   x"90",   x"8A",   x"0E",   x"41",   x"C5", 
  x"75",   x"F1",   x"BE",   x"3A",   x"20",   x"A4",   x"EB",   x"6F", 
  x"48",   x"CC",   x"83",   x"07",   x"1D",   x"99",   x"D6",   x"52", 
  x"E2",   x"66",   x"29",   x"AD",   x"B7",   x"33",   x"7C",   x"F8", 
  x"2B",   x"AF",   x"E0",   x"64",   x"7E",   x"FA",   x"B5",   x"31", 
  x"81",   x"05",   x"4A",   x"CE",   x"D4",   x"50",   x"1F",   x"9B", 
  x"BC",   x"38",   x"77",   x"F3",   x"E9",   x"6D",   x"22",   x"A6", 
  x"16",   x"92",   x"DD",   x"59",   x"43",   x"C7",   x"88",   x"0C", 
  x"C6",   x"42",   x"0D",   x"89",   x"93",   x"17",   x"58",   x"DC", 
  x"6C",   x"E8",   x"A7",   x"23",   x"39",   x"BD",   x"F2",   x"76", 
  x"51",   x"D5",   x"9A",   x"1E",   x"04",   x"80",   x"CF",   x"4B", 
  x"FB",   x"7F",   x"30",   x"B4",   x"AE",   x"2A",   x"65",   x"E1", 
  x"00",   x"85",   x"C9",   x"4C",   x"51",   x"D4",   x"98",   x"1D", 
  x"A2",   x"27",   x"6B",   x"EE",   x"F3",   x"76",   x"3A",   x"BF", 
  x"87",   x"02",   x"4E",   x"CB",   x"D6",   x"53",   x"1F",   x"9A", 
  x"25",   x"A0",   x"EC",   x"69",   x"74",   x"F1",   x"BD",   x"38", 
  x"CD",   x"48",   x"04",   x"81",   x"9C",   x"19",   x"55",   x"D0", 
  x"6F",   x"EA",   x"A6",   x"23",   x"3E",   x"BB",   x"F7",   x"72", 
  x"4A",   x"CF",   x"83",   x"06",   x"1B",   x"9E",   x"D2",   x"57", 
  x"E8",   x"6D",   x"21",   x"A4",   x"B9",   x"3C",   x"70",   x"F5", 
  x"59",   x"DC",   x"90",   x"15",   x"08",   x"8D",   x"C1",   x"44", 
  x"FB",   x"7E",   x"32",   x"B7",   x"AA",   x"2F",   x"63",   x"E6", 
  x"DE",   x"5B",   x"17",   x"92",   x"8F",   x"0A",   x"46",   x"C3", 
  x"7C",   x"F9",   x"B5",   x"30",   x"2D",   x"A8",   x"E4",   x"61", 
  x"94",   x"11",   x"5D",   x"D8",   x"C5",   x"40",   x"0C",   x"89", 
  x"36",   x"B3",   x"FF",   x"7A",   x"67",   x"E2",   x"AE",   x"2B", 
  x"13",   x"96",   x"DA",   x"5F",   x"42",   x"C7",   x"8B",   x"0E", 
  x"B1",   x"34",   x"78",   x"FD",   x"E0",   x"65",   x"29",   x"AC", 
  x"B2",   x"37",   x"7B",   x"FE",   x"E3",   x"66",   x"2A",   x"AF", 
  x"10",   x"95",   x"D9",   x"5C",   x"41",   x"C4",   x"88",   x"0D", 
  x"35",   x"B0",   x"FC",   x"79",   x"64",   x"E1",   x"AD",   x"28", 
  x"97",   x"12",   x"5E",   x"DB",   x"C6",   x"43",   x"0F",   x"8A", 
  x"7F",   x"FA",   x"B6",   x"33",   x"2E",   x"AB",   x"E7",   x"62", 
  x"DD",   x"58",   x"14",   x"91",   x"8C",   x"09",   x"45",   x"C0", 
  x"F8",   x"7D",   x"31",   x"B4",   x"A9",   x"2C",   x"60",   x"E5", 
  x"5A",   x"DF",   x"93",   x"16",   x"0B",   x"8E",   x"C2",   x"47", 
  x"EB",   x"6E",   x"22",   x"A7",   x"BA",   x"3F",   x"73",   x"F6", 
  x"49",   x"CC",   x"80",   x"05",   x"18",   x"9D",   x"D1",   x"54", 
  x"6C",   x"E9",   x"A5",   x"20",   x"3D",   x"B8",   x"F4",   x"71", 
  x"CE",   x"4B",   x"07",   x"82",   x"9F",   x"1A",   x"56",   x"D3", 
  x"26",   x"A3",   x"EF",   x"6A",   x"77",   x"F2",   x"BE",   x"3B", 
  x"84",   x"01",   x"4D",   x"C8",   x"D5",   x"50",   x"1C",   x"99", 
  x"A1",   x"24",   x"68",   x"ED",   x"F0",   x"75",   x"39",   x"BC", 
  x"03",   x"86",   x"CA",   x"4F",   x"52",   x"D7",   x"9B",   x"1E", 
  x"00",   x"86",   x"CF",   x"49",   x"5D",   x"DB",   x"92",   x"14", 
  x"BA",   x"3C",   x"75",   x"F3",   x"E7",   x"61",   x"28",   x"AE", 
  x"B7",   x"31",   x"78",   x"FE",   x"EA",   x"6C",   x"25",   x"A3", 
  x"0D",   x"8B",   x"C2",   x"44",   x"50",   x"D6",   x"9F",   x"19", 
  x"AD",   x"2B",   x"62",   x"E4",   x"F0",   x"76",   x"3F",   x"B9", 
  x"17",   x"91",   x"D8",   x"5E",   x"4A",   x"CC",   x"85",   x"03", 
  x"1A",   x"9C",   x"D5",   x"53",   x"47",   x"C1",   x"88",   x"0E", 
  x"A0",   x"26",   x"6F",   x"E9",   x"FD",   x"7B",   x"32",   x"B4", 
  x"99",   x"1F",   x"56",   x"D0",   x"C4",   x"42",   x"0B",   x"8D", 
  x"23",   x"A5",   x"EC",   x"6A",   x"7E",   x"F8",   x"B1",   x"37", 
  x"2E",   x"A8",   x"E1",   x"67",   x"73",   x"F5",   x"BC",   x"3A", 
  x"94",   x"12",   x"5B",   x"DD",   x"C9",   x"4F",   x"06",   x"80", 
  x"34",   x"B2",   x"FB",   x"7D",   x"69",   x"EF",   x"A6",   x"20", 
  x"8E",   x"08",   x"41",   x"C7",   x"D3",   x"55",   x"1C",   x"9A", 
  x"83",   x"05",   x"4C",   x"CA",   x"DE",   x"58",   x"11",   x"97", 
  x"39",   x"BF",   x"F6",   x"70",   x"64",   x"E2",   x"AB",   x"2D", 
  x"F1",   x"77",   x"3E",   x"B8",   x"AC",   x"2A",   x"63",   x"E5", 
  x"4B",   x"CD",   x"84",   x"02",   x"16",   x"90",   x"D9",   x"5F", 
  x"46",   x"C0",   x"89",   x"0F",   x"1B",   x"9D",   x"D4",   x"52", 
  x"FC",   x"7A",   x"33",   x"B5",   x"A1",   x"27",   x"6E",   x"E8", 
  x"5C",   x"DA",   x"93",   x"15",   x"01",   x"87",   x"CE",   x"48", 
  x"E6",   x"60",   x"29",   x"AF",   x"BB",   x"3D",   x"74",   x"F2", 
  x"EB",   x"6D",   x"24",   x"A2",   x"B6",   x"30",   x"79",   x"FF", 
  x"51",   x"D7",   x"9E",   x"18",   x"0C",   x"8A",   x"C3",   x"45", 
  x"68",   x"EE",   x"A7",   x"21",   x"35",   x"B3",   x"FA",   x"7C", 
  x"D2",   x"54",   x"1D",   x"9B",   x"8F",   x"09",   x"40",   x"C6", 
  x"DF",   x"59",   x"10",   x"96",   x"82",   x"04",   x"4D",   x"CB", 
  x"65",   x"E3",   x"AA",   x"2C",   x"38",   x"BE",   x"F7",   x"71", 
  x"C5",   x"43",   x"0A",   x"8C",   x"98",   x"1E",   x"57",   x"D1", 
  x"7F",   x"F9",   x"B0",   x"36",   x"22",   x"A4",   x"ED",   x"6B", 
  x"72",   x"F4",   x"BD",   x"3B",   x"2F",   x"A9",   x"E0",   x"66", 
  x"C8",   x"4E",   x"07",   x"81",   x"95",   x"13",   x"5A",   x"DC", 
  x"00",   x"87",   x"CD",   x"4A",   x"59",   x"DE",   x"94",   x"13", 
  x"B2",   x"35",   x"7F",   x"F8",   x"EB",   x"6C",   x"26",   x"A1", 
  x"A7",   x"20",   x"6A",   x"ED",   x"FE",   x"79",   x"33",   x"B4", 
  x"15",   x"92",   x"D8",   x"5F",   x"4C",   x"CB",   x"81",   x"06", 
  x"8D",   x"0A",   x"40",   x"C7",   x"D4",   x"53",   x"19",   x"9E", 
  x"3F",   x"B8",   x"F2",   x"75",   x"66",   x"E1",   x"AB",   x"2C", 
  x"2A",   x"AD",   x"E7",   x"60",   x"73",   x"F4",   x"BE",   x"39", 
  x"98",   x"1F",   x"55",   x"D2",   x"C1",   x"46",   x"0C",   x"8B", 
  x"D9",   x"5E",   x"14",   x"93",   x"80",   x"07",   x"4D",   x"CA", 
  x"6B",   x"EC",   x"A6",   x"21",   x"32",   x"B5",   x"FF",   x"78", 
  x"7E",   x"F9",   x"B3",   x"34",   x"27",   x"A0",   x"EA",   x"6D", 
  x"CC",   x"4B",   x"01",   x"86",   x"95",   x"12",   x"58",   x"DF", 
  x"54",   x"D3",   x"99",   x"1E",   x"0D",   x"8A",   x"C0",   x"47", 
  x"E6",   x"61",   x"2B",   x"AC",   x"BF",   x"38",   x"72",   x"F5", 
  x"F3",   x"74",   x"3E",   x"B9",   x"AA",   x"2D",   x"67",   x"E0", 
  x"41",   x"C6",   x"8C",   x"0B",   x"18",   x"9F",   x"D5",   x"52", 
  x"71",   x"F6",   x"BC",   x"3B",   x"28",   x"AF",   x"E5",   x"62", 
  x"C3",   x"44",   x"0E",   x"89",   x"9A",   x"1D",   x"57",   x"D0", 
  x"D6",   x"51",   x"1B",   x"9C",   x"8F",   x"08",   x"42",   x"C5", 
  x"64",   x"E3",   x"A9",   x"2E",   x"3D",   x"BA",   x"F0",   x"77", 
  x"FC",   x"7B",   x"31",   x"B6",   x"A5",   x"22",   x"68",   x"EF", 
  x"4E",   x"C9",   x"83",   x"04",   x"17",   x"90",   x"DA",   x"5D", 
  x"5B",   x"DC",   x"96",   x"11",   x"02",   x"85",   x"CF",   x"48", 
  x"E9",   x"6E",   x"24",   x"A3",   x"B0",   x"37",   x"7D",   x"FA", 
  x"A8",   x"2F",   x"65",   x"E2",   x"F1",   x"76",   x"3C",   x"BB", 
  x"1A",   x"9D",   x"D7",   x"50",   x"43",   x"C4",   x"8E",   x"09", 
  x"0F",   x"88",   x"C2",   x"45",   x"56",   x"D1",   x"9B",   x"1C", 
  x"BD",   x"3A",   x"70",   x"F7",   x"E4",   x"63",   x"29",   x"AE", 
  x"25",   x"A2",   x"E8",   x"6F",   x"7C",   x"FB",   x"B1",   x"36", 
  x"97",   x"10",   x"5A",   x"DD",   x"CE",   x"49",   x"03",   x"84", 
  x"82",   x"05",   x"4F",   x"C8",   x"DB",   x"5C",   x"16",   x"91", 
  x"30",   x"B7",   x"FD",   x"7A",   x"69",   x"EE",   x"A4",   x"23", 
  x"00",   x"88",   x"D3",   x"5B",   x"65",   x"ED",   x"B6",   x"3E", 
  x"CA",   x"42",   x"19",   x"91",   x"AF",   x"27",   x"7C",   x"F4", 
  x"57",   x"DF",   x"84",   x"0C",   x"32",   x"BA",   x"E1",   x"69", 
  x"9D",   x"15",   x"4E",   x"C6",   x"F8",   x"70",   x"2B",   x"A3", 
  x"AE",   x"26",   x"7D",   x"F5",   x"CB",   x"43",   x"18",   x"90", 
  x"64",   x"EC",   x"B7",   x"3F",   x"01",   x"89",   x"D2",   x"5A", 
  x"F9",   x"71",   x"2A",   x"A2",   x"9C",   x"14",   x"4F",   x"C7", 
  x"33",   x"BB",   x"E0",   x"68",   x"56",   x"DE",   x"85",   x"0D", 
  x"9F",   x"17",   x"4C",   x"C4",   x"FA",   x"72",   x"29",   x"A1", 
  x"55",   x"DD",   x"86",   x"0E",   x"30",   x"B8",   x"E3",   x"6B", 
  x"C8",   x"40",   x"1B",   x"93",   x"AD",   x"25",   x"7E",   x"F6", 
  x"02",   x"8A",   x"D1",   x"59",   x"67",   x"EF",   x"B4",   x"3C", 
  x"31",   x"B9",   x"E2",   x"6A",   x"54",   x"DC",   x"87",   x"0F", 
  x"FB",   x"73",   x"28",   x"A0",   x"9E",   x"16",   x"4D",   x"C5", 
  x"66",   x"EE",   x"B5",   x"3D",   x"03",   x"8B",   x"D0",   x"58", 
  x"AC",   x"24",   x"7F",   x"F7",   x"C9",   x"41",   x"1A",   x"92", 
  x"FD",   x"75",   x"2E",   x"A6",   x"98",   x"10",   x"4B",   x"C3", 
  x"37",   x"BF",   x"E4",   x"6C",   x"52",   x"DA",   x"81",   x"09", 
  x"AA",   x"22",   x"79",   x"F1",   x"CF",   x"47",   x"1C",   x"94", 
  x"60",   x"E8",   x"B3",   x"3B",   x"05",   x"8D",   x"D6",   x"5E", 
  x"53",   x"DB",   x"80",   x"08",   x"36",   x"BE",   x"E5",   x"6D", 
  x"99",   x"11",   x"4A",   x"C2",   x"FC",   x"74",   x"2F",   x"A7", 
  x"04",   x"8C",   x"D7",   x"5F",   x"61",   x"E9",   x"B2",   x"3A", 
  x"CE",   x"46",   x"1D",   x"95",   x"AB",   x"23",   x"78",   x"F0", 
  x"62",   x"EA",   x"B1",   x"39",   x"07",   x"8F",   x"D4",   x"5C", 
  x"A8",   x"20",   x"7B",   x"F3",   x"CD",   x"45",   x"1E",   x"96", 
  x"35",   x"BD",   x"E6",   x"6E",   x"50",   x"D8",   x"83",   x"0B", 
  x"FF",   x"77",   x"2C",   x"A4",   x"9A",   x"12",   x"49",   x"C1", 
  x"CC",   x"44",   x"1F",   x"97",   x"A9",   x"21",   x"7A",   x"F2", 
  x"06",   x"8E",   x"D5",   x"5D",   x"63",   x"EB",   x"B0",   x"38", 
  x"9B",   x"13",   x"48",   x"C0",   x"FE",   x"76",   x"2D",   x"A5", 
  x"51",   x"D9",   x"82",   x"0A",   x"34",   x"BC",   x"E7",   x"6F", 
  x"00",   x"89",   x"D1",   x"58",   x"61",   x"E8",   x"B0",   x"39", 
  x"C2",   x"4B",   x"13",   x"9A",   x"A3",   x"2A",   x"72",   x"FB", 
  x"47",   x"CE",   x"96",   x"1F",   x"26",   x"AF",   x"F7",   x"7E", 
  x"85",   x"0C",   x"54",   x"DD",   x"E4",   x"6D",   x"35",   x"BC", 
  x"8E",   x"07",   x"5F",   x"D6",   x"EF",   x"66",   x"3E",   x"B7", 
  x"4C",   x"C5",   x"9D",   x"14",   x"2D",   x"A4",   x"FC",   x"75", 
  x"C9",   x"40",   x"18",   x"91",   x"A8",   x"21",   x"79",   x"F0", 
  x"0B",   x"82",   x"DA",   x"53",   x"6A",   x"E3",   x"BB",   x"32", 
  x"DF",   x"56",   x"0E",   x"87",   x"BE",   x"37",   x"6F",   x"E6", 
  x"1D",   x"94",   x"CC",   x"45",   x"7C",   x"F5",   x"AD",   x"24", 
  x"98",   x"11",   x"49",   x"C0",   x"F9",   x"70",   x"28",   x"A1", 
  x"5A",   x"D3",   x"8B",   x"02",   x"3B",   x"B2",   x"EA",   x"63", 
  x"51",   x"D8",   x"80",   x"09",   x"30",   x"B9",   x"E1",   x"68", 
  x"93",   x"1A",   x"42",   x"CB",   x"F2",   x"7B",   x"23",   x"AA", 
  x"16",   x"9F",   x"C7",   x"4E",   x"77",   x"FE",   x"A6",   x"2F", 
  x"D4",   x"5D",   x"05",   x"8C",   x"B5",   x"3C",   x"64",   x"ED", 
  x"7D",   x"F4",   x"AC",   x"25",   x"1C",   x"95",   x"CD",   x"44", 
  x"BF",   x"36",   x"6E",   x"E7",   x"DE",   x"57",   x"0F",   x"86", 
  x"3A",   x"B3",   x"EB",   x"62",   x"5B",   x"D2",   x"8A",   x"03", 
  x"F8",   x"71",   x"29",   x"A0",   x"99",   x"10",   x"48",   x"C1", 
  x"F3",   x"7A",   x"22",   x"AB",   x"92",   x"1B",   x"43",   x"CA", 
  x"31",   x"B8",   x"E0",   x"69",   x"50",   x"D9",   x"81",   x"08", 
  x"B4",   x"3D",   x"65",   x"EC",   x"D5",   x"5C",   x"04",   x"8D", 
  x"76",   x"FF",   x"A7",   x"2E",   x"17",   x"9E",   x"C6",   x"4F", 
  x"A2",   x"2B",   x"73",   x"FA",   x"C3",   x"4A",   x"12",   x"9B", 
  x"60",   x"E9",   x"B1",   x"38",   x"01",   x"88",   x"D0",   x"59", 
  x"E5",   x"6C",   x"34",   x"BD",   x"84",   x"0D",   x"55",   x"DC", 
  x"27",   x"AE",   x"F6",   x"7F",   x"46",   x"CF",   x"97",   x"1E", 
  x"2C",   x"A5",   x"FD",   x"74",   x"4D",   x"C4",   x"9C",   x"15", 
  x"EE",   x"67",   x"3F",   x"B6",   x"8F",   x"06",   x"5E",   x"D7", 
  x"6B",   x"E2",   x"BA",   x"33",   x"0A",   x"83",   x"DB",   x"52", 
  x"A9",   x"20",   x"78",   x"F1",   x"C8",   x"41",   x"19",   x"90", 
  x"00",   x"8A",   x"D7",   x"5D",   x"6D",   x"E7",   x"BA",   x"30", 
  x"DA",   x"50",   x"0D",   x"87",   x"B7",   x"3D",   x"60",   x"EA", 
  x"77",   x"FD",   x"A0",   x"2A",   x"1A",   x"90",   x"CD",   x"47", 
  x"AD",   x"27",   x"7A",   x"F0",   x"C0",   x"4A",   x"17",   x"9D", 
  x"EE",   x"64",   x"39",   x"B3",   x"83",   x"09",   x"54",   x"DE", 
  x"34",   x"BE",   x"E3",   x"69",   x"59",   x"D3",   x"8E",   x"04", 
  x"99",   x"13",   x"4E",   x"C4",   x"F4",   x"7E",   x"23",   x"A9", 
  x"43",   x"C9",   x"94",   x"1E",   x"2E",   x"A4",   x"F9",   x"73", 
  x"1F",   x"95",   x"C8",   x"42",   x"72",   x"F8",   x"A5",   x"2F", 
  x"C5",   x"4F",   x"12",   x"98",   x"A8",   x"22",   x"7F",   x"F5", 
  x"68",   x"E2",   x"BF",   x"35",   x"05",   x"8F",   x"D2",   x"58", 
  x"B2",   x"38",   x"65",   x"EF",   x"DF",   x"55",   x"08",   x"82", 
  x"F1",   x"7B",   x"26",   x"AC",   x"9C",   x"16",   x"4B",   x"C1", 
  x"2B",   x"A1",   x"FC",   x"76",   x"46",   x"CC",   x"91",   x"1B", 
  x"86",   x"0C",   x"51",   x"DB",   x"EB",   x"61",   x"3C",   x"B6", 
  x"5C",   x"D6",   x"8B",   x"01",   x"31",   x"BB",   x"E6",   x"6C", 
  x"3E",   x"B4",   x"E9",   x"63",   x"53",   x"D9",   x"84",   x"0E", 
  x"E4",   x"6E",   x"33",   x"B9",   x"89",   x"03",   x"5E",   x"D4", 
  x"49",   x"C3",   x"9E",   x"14",   x"24",   x"AE",   x"F3",   x"79", 
  x"93",   x"19",   x"44",   x"CE",   x"FE",   x"74",   x"29",   x"A3", 
  x"D0",   x"5A",   x"07",   x"8D",   x"BD",   x"37",   x"6A",   x"E0", 
  x"0A",   x"80",   x"DD",   x"57",   x"67",   x"ED",   x"B0",   x"3A", 
  x"A7",   x"2D",   x"70",   x"FA",   x"CA",   x"40",   x"1D",   x"97", 
  x"7D",   x"F7",   x"AA",   x"20",   x"10",   x"9A",   x"C7",   x"4D", 
  x"21",   x"AB",   x"F6",   x"7C",   x"4C",   x"C6",   x"9B",   x"11", 
  x"FB",   x"71",   x"2C",   x"A6",   x"96",   x"1C",   x"41",   x"CB", 
  x"56",   x"DC",   x"81",   x"0B",   x"3B",   x"B1",   x"EC",   x"66", 
  x"8C",   x"06",   x"5B",   x"D1",   x"E1",   x"6B",   x"36",   x"BC", 
  x"CF",   x"45",   x"18",   x"92",   x"A2",   x"28",   x"75",   x"FF", 
  x"15",   x"9F",   x"C2",   x"48",   x"78",   x"F2",   x"AF",   x"25", 
  x"B8",   x"32",   x"6F",   x"E5",   x"D5",   x"5F",   x"02",   x"88", 
  x"62",   x"E8",   x"B5",   x"3F",   x"0F",   x"85",   x"D8",   x"52", 
  x"00",   x"8B",   x"D5",   x"5E",   x"69",   x"E2",   x"BC",   x"37", 
  x"D2",   x"59",   x"07",   x"8C",   x"BB",   x"30",   x"6E",   x"E5", 
  x"67",   x"EC",   x"B2",   x"39",   x"0E",   x"85",   x"DB",   x"50", 
  x"B5",   x"3E",   x"60",   x"EB",   x"DC",   x"57",   x"09",   x"82", 
  x"CE",   x"45",   x"1B",   x"90",   x"A7",   x"2C",   x"72",   x"F9", 
  x"1C",   x"97",   x"C9",   x"42",   x"75",   x"FE",   x"A0",   x"2B", 
  x"A9",   x"22",   x"7C",   x"F7",   x"C0",   x"4B",   x"15",   x"9E", 
  x"7B",   x"F0",   x"AE",   x"25",   x"12",   x"99",   x"C7",   x"4C", 
  x"5F",   x"D4",   x"8A",   x"01",   x"36",   x"BD",   x"E3",   x"68", 
  x"8D",   x"06",   x"58",   x"D3",   x"E4",   x"6F",   x"31",   x"BA", 
  x"38",   x"B3",   x"ED",   x"66",   x"51",   x"DA",   x"84",   x"0F", 
  x"EA",   x"61",   x"3F",   x"B4",   x"83",   x"08",   x"56",   x"DD", 
  x"91",   x"1A",   x"44",   x"CF",   x"F8",   x"73",   x"2D",   x"A6", 
  x"43",   x"C8",   x"96",   x"1D",   x"2A",   x"A1",   x"FF",   x"74", 
  x"F6",   x"7D",   x"23",   x"A8",   x"9F",   x"14",   x"4A",   x"C1", 
  x"24",   x"AF",   x"F1",   x"7A",   x"4D",   x"C6",   x"98",   x"13", 
  x"BE",   x"35",   x"6B",   x"E0",   x"D7",   x"5C",   x"02",   x"89", 
  x"6C",   x"E7",   x"B9",   x"32",   x"05",   x"8E",   x"D0",   x"5B", 
  x"D9",   x"52",   x"0C",   x"87",   x"B0",   x"3B",   x"65",   x"EE", 
  x"0B",   x"80",   x"DE",   x"55",   x"62",   x"E9",   x"B7",   x"3C", 
  x"70",   x"FB",   x"A5",   x"2E",   x"19",   x"92",   x"CC",   x"47", 
  x"A2",   x"29",   x"77",   x"FC",   x"CB",   x"40",   x"1E",   x"95", 
  x"17",   x"9C",   x"C2",   x"49",   x"7E",   x"F5",   x"AB",   x"20", 
  x"C5",   x"4E",   x"10",   x"9B",   x"AC",   x"27",   x"79",   x"F2", 
  x"E1",   x"6A",   x"34",   x"BF",   x"88",   x"03",   x"5D",   x"D6", 
  x"33",   x"B8",   x"E6",   x"6D",   x"5A",   x"D1",   x"8F",   x"04", 
  x"86",   x"0D",   x"53",   x"D8",   x"EF",   x"64",   x"3A",   x"B1", 
  x"54",   x"DF",   x"81",   x"0A",   x"3D",   x"B6",   x"E8",   x"63", 
  x"2F",   x"A4",   x"FA",   x"71",   x"46",   x"CD",   x"93",   x"18", 
  x"FD",   x"76",   x"28",   x"A3",   x"94",   x"1F",   x"41",   x"CA", 
  x"48",   x"C3",   x"9D",   x"16",   x"21",   x"AA",   x"F4",   x"7F", 
  x"9A",   x"11",   x"4F",   x"C4",   x"F3",   x"78",   x"26",   x"AD", 
  x"00",   x"8C",   x"DB",   x"57",   x"75",   x"F9",   x"AE",   x"22", 
  x"EA",   x"66",   x"31",   x"BD",   x"9F",   x"13",   x"44",   x"C8", 
  x"17",   x"9B",   x"CC",   x"40",   x"62",   x"EE",   x"B9",   x"35", 
  x"FD",   x"71",   x"26",   x"AA",   x"88",   x"04",   x"53",   x"DF", 
  x"2E",   x"A2",   x"F5",   x"79",   x"5B",   x"D7",   x"80",   x"0C", 
  x"C4",   x"48",   x"1F",   x"93",   x"B1",   x"3D",   x"6A",   x"E6", 
  x"39",   x"B5",   x"E2",   x"6E",   x"4C",   x"C0",   x"97",   x"1B", 
  x"D3",   x"5F",   x"08",   x"84",   x"A6",   x"2A",   x"7D",   x"F1", 
  x"5C",   x"D0",   x"87",   x"0B",   x"29",   x"A5",   x"F2",   x"7E", 
  x"B6",   x"3A",   x"6D",   x"E1",   x"C3",   x"4F",   x"18",   x"94", 
  x"4B",   x"C7",   x"90",   x"1C",   x"3E",   x"B2",   x"E5",   x"69", 
  x"A1",   x"2D",   x"7A",   x"F6",   x"D4",   x"58",   x"0F",   x"83", 
  x"72",   x"FE",   x"A9",   x"25",   x"07",   x"8B",   x"DC",   x"50", 
  x"98",   x"14",   x"43",   x"CF",   x"ED",   x"61",   x"36",   x"BA", 
  x"65",   x"E9",   x"BE",   x"32",   x"10",   x"9C",   x"CB",   x"47", 
  x"8F",   x"03",   x"54",   x"D8",   x"FA",   x"76",   x"21",   x"AD", 
  x"B8",   x"34",   x"63",   x"EF",   x"CD",   x"41",   x"16",   x"9A", 
  x"52",   x"DE",   x"89",   x"05",   x"27",   x"AB",   x"FC",   x"70", 
  x"AF",   x"23",   x"74",   x"F8",   x"DA",   x"56",   x"01",   x"8D", 
  x"45",   x"C9",   x"9E",   x"12",   x"30",   x"BC",   x"EB",   x"67", 
  x"96",   x"1A",   x"4D",   x"C1",   x"E3",   x"6F",   x"38",   x"B4", 
  x"7C",   x"F0",   x"A7",   x"2B",   x"09",   x"85",   x"D2",   x"5E", 
  x"81",   x"0D",   x"5A",   x"D6",   x"F4",   x"78",   x"2F",   x"A3", 
  x"6B",   x"E7",   x"B0",   x"3C",   x"1E",   x"92",   x"C5",   x"49", 
  x"E4",   x"68",   x"3F",   x"B3",   x"91",   x"1D",   x"4A",   x"C6", 
  x"0E",   x"82",   x"D5",   x"59",   x"7B",   x"F7",   x"A0",   x"2C", 
  x"F3",   x"7F",   x"28",   x"A4",   x"86",   x"0A",   x"5D",   x"D1", 
  x"19",   x"95",   x"C2",   x"4E",   x"6C",   x"E0",   x"B7",   x"3B", 
  x"CA",   x"46",   x"11",   x"9D",   x"BF",   x"33",   x"64",   x"E8", 
  x"20",   x"AC",   x"FB",   x"77",   x"55",   x"D9",   x"8E",   x"02", 
  x"DD",   x"51",   x"06",   x"8A",   x"A8",   x"24",   x"73",   x"FF", 
  x"37",   x"BB",   x"EC",   x"60",   x"42",   x"CE",   x"99",   x"15", 
  x"00",   x"8D",   x"D9",   x"54",   x"71",   x"FC",   x"A8",   x"25", 
  x"E2",   x"6F",   x"3B",   x"B6",   x"93",   x"1E",   x"4A",   x"C7", 
  x"07",   x"8A",   x"DE",   x"53",   x"76",   x"FB",   x"AF",   x"22", 
  x"E5",   x"68",   x"3C",   x"B1",   x"94",   x"19",   x"4D",   x"C0", 
  x"0E",   x"83",   x"D7",   x"5A",   x"7F",   x"F2",   x"A6",   x"2B", 
  x"EC",   x"61",   x"35",   x"B8",   x"9D",   x"10",   x"44",   x"C9", 
  x"09",   x"84",   x"D0",   x"5D",   x"78",   x"F5",   x"A1",   x"2C", 
  x"EB",   x"66",   x"32",   x"BF",   x"9A",   x"17",   x"43",   x"CE", 
  x"1C",   x"91",   x"C5",   x"48",   x"6D",   x"E0",   x"B4",   x"39", 
  x"FE",   x"73",   x"27",   x"AA",   x"8F",   x"02",   x"56",   x"DB", 
  x"1B",   x"96",   x"C2",   x"4F",   x"6A",   x"E7",   x"B3",   x"3E", 
  x"F9",   x"74",   x"20",   x"AD",   x"88",   x"05",   x"51",   x"DC", 
  x"12",   x"9F",   x"CB",   x"46",   x"63",   x"EE",   x"BA",   x"37", 
  x"F0",   x"7D",   x"29",   x"A4",   x"81",   x"0C",   x"58",   x"D5", 
  x"15",   x"98",   x"CC",   x"41",   x"64",   x"E9",   x"BD",   x"30", 
  x"F7",   x"7A",   x"2E",   x"A3",   x"86",   x"0B",   x"5F",   x"D2", 
  x"38",   x"B5",   x"E1",   x"6C",   x"49",   x"C4",   x"90",   x"1D", 
  x"DA",   x"57",   x"03",   x"8E",   x"AB",   x"26",   x"72",   x"FF", 
  x"3F",   x"B2",   x"E6",   x"6B",   x"4E",   x"C3",   x"97",   x"1A", 
  x"DD",   x"50",   x"04",   x"89",   x"AC",   x"21",   x"75",   x"F8", 
  x"36",   x"BB",   x"EF",   x"62",   x"47",   x"CA",   x"9E",   x"13", 
  x"D4",   x"59",   x"0D",   x"80",   x"A5",   x"28",   x"7C",   x"F1", 
  x"31",   x"BC",   x"E8",   x"65",   x"40",   x"CD",   x"99",   x"14", 
  x"D3",   x"5E",   x"0A",   x"87",   x"A2",   x"2F",   x"7B",   x"F6", 
  x"24",   x"A9",   x"FD",   x"70",   x"55",   x"D8",   x"8C",   x"01", 
  x"C6",   x"4B",   x"1F",   x"92",   x"B7",   x"3A",   x"6E",   x"E3", 
  x"23",   x"AE",   x"FA",   x"77",   x"52",   x"DF",   x"8B",   x"06", 
  x"C1",   x"4C",   x"18",   x"95",   x"B0",   x"3D",   x"69",   x"E4", 
  x"2A",   x"A7",   x"F3",   x"7E",   x"5B",   x"D6",   x"82",   x"0F", 
  x"C8",   x"45",   x"11",   x"9C",   x"B9",   x"34",   x"60",   x"ED", 
  x"2D",   x"A0",   x"F4",   x"79",   x"5C",   x"D1",   x"85",   x"08", 
  x"CF",   x"42",   x"16",   x"9B",   x"BE",   x"33",   x"67",   x"EA", 
  x"00",   x"8E",   x"DF",   x"51",   x"7D",   x"F3",   x"A2",   x"2C", 
  x"FA",   x"74",   x"25",   x"AB",   x"87",   x"09",   x"58",   x"D6", 
  x"37",   x"B9",   x"E8",   x"66",   x"4A",   x"C4",   x"95",   x"1B", 
  x"CD",   x"43",   x"12",   x"9C",   x"B0",   x"3E",   x"6F",   x"E1", 
  x"6E",   x"E0",   x"B1",   x"3F",   x"13",   x"9D",   x"CC",   x"42", 
  x"94",   x"1A",   x"4B",   x"C5",   x"E9",   x"67",   x"36",   x"B8", 
  x"59",   x"D7",   x"86",   x"08",   x"24",   x"AA",   x"FB",   x"75", 
  x"A3",   x"2D",   x"7C",   x"F2",   x"DE",   x"50",   x"01",   x"8F", 
  x"DC",   x"52",   x"03",   x"8D",   x"A1",   x"2F",   x"7E",   x"F0", 
  x"26",   x"A8",   x"F9",   x"77",   x"5B",   x"D5",   x"84",   x"0A", 
  x"EB",   x"65",   x"34",   x"BA",   x"96",   x"18",   x"49",   x"C7", 
  x"11",   x"9F",   x"CE",   x"40",   x"6C",   x"E2",   x"B3",   x"3D", 
  x"B2",   x"3C",   x"6D",   x"E3",   x"CF",   x"41",   x"10",   x"9E", 
  x"48",   x"C6",   x"97",   x"19",   x"35",   x"BB",   x"EA",   x"64", 
  x"85",   x"0B",   x"5A",   x"D4",   x"F8",   x"76",   x"27",   x"A9", 
  x"7F",   x"F1",   x"A0",   x"2E",   x"02",   x"8C",   x"DD",   x"53", 
  x"7B",   x"F5",   x"A4",   x"2A",   x"06",   x"88",   x"D9",   x"57", 
  x"81",   x"0F",   x"5E",   x"D0",   x"FC",   x"72",   x"23",   x"AD", 
  x"4C",   x"C2",   x"93",   x"1D",   x"31",   x"BF",   x"EE",   x"60", 
  x"B6",   x"38",   x"69",   x"E7",   x"CB",   x"45",   x"14",   x"9A", 
  x"15",   x"9B",   x"CA",   x"44",   x"68",   x"E6",   x"B7",   x"39", 
  x"EF",   x"61",   x"30",   x"BE",   x"92",   x"1C",   x"4D",   x"C3", 
  x"22",   x"AC",   x"FD",   x"73",   x"5F",   x"D1",   x"80",   x"0E", 
  x"D8",   x"56",   x"07",   x"89",   x"A5",   x"2B",   x"7A",   x"F4", 
  x"A7",   x"29",   x"78",   x"F6",   x"DA",   x"54",   x"05",   x"8B", 
  x"5D",   x"D3",   x"82",   x"0C",   x"20",   x"AE",   x"FF",   x"71", 
  x"90",   x"1E",   x"4F",   x"C1",   x"ED",   x"63",   x"32",   x"BC", 
  x"6A",   x"E4",   x"B5",   x"3B",   x"17",   x"99",   x"C8",   x"46", 
  x"C9",   x"47",   x"16",   x"98",   x"B4",   x"3A",   x"6B",   x"E5", 
  x"33",   x"BD",   x"EC",   x"62",   x"4E",   x"C0",   x"91",   x"1F", 
  x"FE",   x"70",   x"21",   x"AF",   x"83",   x"0D",   x"5C",   x"D2", 
  x"04",   x"8A",   x"DB",   x"55",   x"79",   x"F7",   x"A6",   x"28", 
  x"00",   x"8F",   x"DD",   x"52",   x"79",   x"F6",   x"A4",   x"2B", 
  x"F2",   x"7D",   x"2F",   x"A0",   x"8B",   x"04",   x"56",   x"D9", 
  x"27",   x"A8",   x"FA",   x"75",   x"5E",   x"D1",   x"83",   x"0C", 
  x"D5",   x"5A",   x"08",   x"87",   x"AC",   x"23",   x"71",   x"FE", 
  x"4E",   x"C1",   x"93",   x"1C",   x"37",   x"B8",   x"EA",   x"65", 
  x"BC",   x"33",   x"61",   x"EE",   x"C5",   x"4A",   x"18",   x"97", 
  x"69",   x"E6",   x"B4",   x"3B",   x"10",   x"9F",   x"CD",   x"42", 
  x"9B",   x"14",   x"46",   x"C9",   x"E2",   x"6D",   x"3F",   x"B0", 
  x"9C",   x"13",   x"41",   x"CE",   x"E5",   x"6A",   x"38",   x"B7", 
  x"6E",   x"E1",   x"B3",   x"3C",   x"17",   x"98",   x"CA",   x"45", 
  x"BB",   x"34",   x"66",   x"E9",   x"C2",   x"4D",   x"1F",   x"90", 
  x"49",   x"C6",   x"94",   x"1B",   x"30",   x"BF",   x"ED",   x"62", 
  x"D2",   x"5D",   x"0F",   x"80",   x"AB",   x"24",   x"76",   x"F9", 
  x"20",   x"AF",   x"FD",   x"72",   x"59",   x"D6",   x"84",   x"0B", 
  x"F5",   x"7A",   x"28",   x"A7",   x"8C",   x"03",   x"51",   x"DE", 
  x"07",   x"88",   x"DA",   x"55",   x"7E",   x"F1",   x"A3",   x"2C", 
  x"FB",   x"74",   x"26",   x"A9",   x"82",   x"0D",   x"5F",   x"D0", 
  x"09",   x"86",   x"D4",   x"5B",   x"70",   x"FF",   x"AD",   x"22", 
  x"DC",   x"53",   x"01",   x"8E",   x"A5",   x"2A",   x"78",   x"F7", 
  x"2E",   x"A1",   x"F3",   x"7C",   x"57",   x"D8",   x"8A",   x"05", 
  x"B5",   x"3A",   x"68",   x"E7",   x"CC",   x"43",   x"11",   x"9E", 
  x"47",   x"C8",   x"9A",   x"15",   x"3E",   x"B1",   x"E3",   x"6C", 
  x"92",   x"1D",   x"4F",   x"C0",   x"EB",   x"64",   x"36",   x"B9", 
  x"60",   x"EF",   x"BD",   x"32",   x"19",   x"96",   x"C4",   x"4B", 
  x"67",   x"E8",   x"BA",   x"35",   x"1E",   x"91",   x"C3",   x"4C", 
  x"95",   x"1A",   x"48",   x"C7",   x"EC",   x"63",   x"31",   x"BE", 
  x"40",   x"CF",   x"9D",   x"12",   x"39",   x"B6",   x"E4",   x"6B", 
  x"B2",   x"3D",   x"6F",   x"E0",   x"CB",   x"44",   x"16",   x"99", 
  x"29",   x"A6",   x"F4",   x"7B",   x"50",   x"DF",   x"8D",   x"02", 
  x"DB",   x"54",   x"06",   x"89",   x"A2",   x"2D",   x"7F",   x"F0", 
  x"0E",   x"81",   x"D3",   x"5C",   x"77",   x"F8",   x"AA",   x"25", 
  x"FC",   x"73",   x"21",   x"AE",   x"85",   x"0A",   x"58",   x"D7", 
  x"00",   x"90",   x"E3",   x"73",   x"05",   x"95",   x"E6",   x"76", 
  x"0A",   x"9A",   x"E9",   x"79",   x"0F",   x"9F",   x"EC",   x"7C", 
  x"14",   x"84",   x"F7",   x"67",   x"11",   x"81",   x"F2",   x"62", 
  x"1E",   x"8E",   x"FD",   x"6D",   x"1B",   x"8B",   x"F8",   x"68", 
  x"28",   x"B8",   x"CB",   x"5B",   x"2D",   x"BD",   x"CE",   x"5E", 
  x"22",   x"B2",   x"C1",   x"51",   x"27",   x"B7",   x"C4",   x"54", 
  x"3C",   x"AC",   x"DF",   x"4F",   x"39",   x"A9",   x"DA",   x"4A", 
  x"36",   x"A6",   x"D5",   x"45",   x"33",   x"A3",   x"D0",   x"40", 
  x"50",   x"C0",   x"B3",   x"23",   x"55",   x"C5",   x"B6",   x"26", 
  x"5A",   x"CA",   x"B9",   x"29",   x"5F",   x"CF",   x"BC",   x"2C", 
  x"44",   x"D4",   x"A7",   x"37",   x"41",   x"D1",   x"A2",   x"32", 
  x"4E",   x"DE",   x"AD",   x"3D",   x"4B",   x"DB",   x"A8",   x"38", 
  x"78",   x"E8",   x"9B",   x"0B",   x"7D",   x"ED",   x"9E",   x"0E", 
  x"72",   x"E2",   x"91",   x"01",   x"77",   x"E7",   x"94",   x"04", 
  x"6C",   x"FC",   x"8F",   x"1F",   x"69",   x"F9",   x"8A",   x"1A", 
  x"66",   x"F6",   x"85",   x"15",   x"63",   x"F3",   x"80",   x"10", 
  x"A0",   x"30",   x"43",   x"D3",   x"A5",   x"35",   x"46",   x"D6", 
  x"AA",   x"3A",   x"49",   x"D9",   x"AF",   x"3F",   x"4C",   x"DC", 
  x"B4",   x"24",   x"57",   x"C7",   x"B1",   x"21",   x"52",   x"C2", 
  x"BE",   x"2E",   x"5D",   x"CD",   x"BB",   x"2B",   x"58",   x"C8", 
  x"88",   x"18",   x"6B",   x"FB",   x"8D",   x"1D",   x"6E",   x"FE", 
  x"82",   x"12",   x"61",   x"F1",   x"87",   x"17",   x"64",   x"F4", 
  x"9C",   x"0C",   x"7F",   x"EF",   x"99",   x"09",   x"7A",   x"EA", 
  x"96",   x"06",   x"75",   x"E5",   x"93",   x"03",   x"70",   x"E0", 
  x"F0",   x"60",   x"13",   x"83",   x"F5",   x"65",   x"16",   x"86", 
  x"FA",   x"6A",   x"19",   x"89",   x"FF",   x"6F",   x"1C",   x"8C", 
  x"E4",   x"74",   x"07",   x"97",   x"E1",   x"71",   x"02",   x"92", 
  x"EE",   x"7E",   x"0D",   x"9D",   x"EB",   x"7B",   x"08",   x"98", 
  x"D8",   x"48",   x"3B",   x"AB",   x"DD",   x"4D",   x"3E",   x"AE", 
  x"D2",   x"42",   x"31",   x"A1",   x"D7",   x"47",   x"34",   x"A4", 
  x"CC",   x"5C",   x"2F",   x"BF",   x"C9",   x"59",   x"2A",   x"BA", 
  x"C6",   x"56",   x"25",   x"B5",   x"C3",   x"53",   x"20",   x"B0", 
  x"00",   x"91",   x"E1",   x"70",   x"01",   x"90",   x"E0",   x"71", 
  x"02",   x"93",   x"E3",   x"72",   x"03",   x"92",   x"E2",   x"73", 
  x"04",   x"95",   x"E5",   x"74",   x"05",   x"94",   x"E4",   x"75", 
  x"06",   x"97",   x"E7",   x"76",   x"07",   x"96",   x"E6",   x"77", 
  x"08",   x"99",   x"E9",   x"78",   x"09",   x"98",   x"E8",   x"79", 
  x"0A",   x"9B",   x"EB",   x"7A",   x"0B",   x"9A",   x"EA",   x"7B", 
  x"0C",   x"9D",   x"ED",   x"7C",   x"0D",   x"9C",   x"EC",   x"7D", 
  x"0E",   x"9F",   x"EF",   x"7E",   x"0F",   x"9E",   x"EE",   x"7F", 
  x"10",   x"81",   x"F1",   x"60",   x"11",   x"80",   x"F0",   x"61", 
  x"12",   x"83",   x"F3",   x"62",   x"13",   x"82",   x"F2",   x"63", 
  x"14",   x"85",   x"F5",   x"64",   x"15",   x"84",   x"F4",   x"65", 
  x"16",   x"87",   x"F7",   x"66",   x"17",   x"86",   x"F6",   x"67", 
  x"18",   x"89",   x"F9",   x"68",   x"19",   x"88",   x"F8",   x"69", 
  x"1A",   x"8B",   x"FB",   x"6A",   x"1B",   x"8A",   x"FA",   x"6B", 
  x"1C",   x"8D",   x"FD",   x"6C",   x"1D",   x"8C",   x"FC",   x"6D", 
  x"1E",   x"8F",   x"FF",   x"6E",   x"1F",   x"8E",   x"FE",   x"6F", 
  x"20",   x"B1",   x"C1",   x"50",   x"21",   x"B0",   x"C0",   x"51", 
  x"22",   x"B3",   x"C3",   x"52",   x"23",   x"B2",   x"C2",   x"53", 
  x"24",   x"B5",   x"C5",   x"54",   x"25",   x"B4",   x"C4",   x"55", 
  x"26",   x"B7",   x"C7",   x"56",   x"27",   x"B6",   x"C6",   x"57", 
  x"28",   x"B9",   x"C9",   x"58",   x"29",   x"B8",   x"C8",   x"59", 
  x"2A",   x"BB",   x"CB",   x"5A",   x"2B",   x"BA",   x"CA",   x"5B", 
  x"2C",   x"BD",   x"CD",   x"5C",   x"2D",   x"BC",   x"CC",   x"5D", 
  x"2E",   x"BF",   x"CF",   x"5E",   x"2F",   x"BE",   x"CE",   x"5F", 
  x"30",   x"A1",   x"D1",   x"40",   x"31",   x"A0",   x"D0",   x"41", 
  x"32",   x"A3",   x"D3",   x"42",   x"33",   x"A2",   x"D2",   x"43", 
  x"34",   x"A5",   x"D5",   x"44",   x"35",   x"A4",   x"D4",   x"45", 
  x"36",   x"A7",   x"D7",   x"46",   x"37",   x"A6",   x"D6",   x"47", 
  x"38",   x"A9",   x"D9",   x"48",   x"39",   x"A8",   x"D8",   x"49", 
  x"3A",   x"AB",   x"DB",   x"4A",   x"3B",   x"AA",   x"DA",   x"4B", 
  x"3C",   x"AD",   x"DD",   x"4C",   x"3D",   x"AC",   x"DC",   x"4D", 
  x"3E",   x"AF",   x"DF",   x"4E",   x"3F",   x"AE",   x"DE",   x"4F", 
  x"00",   x"92",   x"E7",   x"75",   x"0D",   x"9F",   x"EA",   x"78", 
  x"1A",   x"88",   x"FD",   x"6F",   x"17",   x"85",   x"F0",   x"62", 
  x"34",   x"A6",   x"D3",   x"41",   x"39",   x"AB",   x"DE",   x"4C", 
  x"2E",   x"BC",   x"C9",   x"5B",   x"23",   x"B1",   x"C4",   x"56", 
  x"68",   x"FA",   x"8F",   x"1D",   x"65",   x"F7",   x"82",   x"10", 
  x"72",   x"E0",   x"95",   x"07",   x"7F",   x"ED",   x"98",   x"0A", 
  x"5C",   x"CE",   x"BB",   x"29",   x"51",   x"C3",   x"B6",   x"24", 
  x"46",   x"D4",   x"A1",   x"33",   x"4B",   x"D9",   x"AC",   x"3E", 
  x"D0",   x"42",   x"37",   x"A5",   x"DD",   x"4F",   x"3A",   x"A8", 
  x"CA",   x"58",   x"2D",   x"BF",   x"C7",   x"55",   x"20",   x"B2", 
  x"E4",   x"76",   x"03",   x"91",   x"E9",   x"7B",   x"0E",   x"9C", 
  x"FE",   x"6C",   x"19",   x"8B",   x"F3",   x"61",   x"14",   x"86", 
  x"B8",   x"2A",   x"5F",   x"CD",   x"B5",   x"27",   x"52",   x"C0", 
  x"A2",   x"30",   x"45",   x"D7",   x"AF",   x"3D",   x"48",   x"DA", 
  x"8C",   x"1E",   x"6B",   x"F9",   x"81",   x"13",   x"66",   x"F4", 
  x"96",   x"04",   x"71",   x"E3",   x"9B",   x"09",   x"7C",   x"EE", 
  x"63",   x"F1",   x"84",   x"16",   x"6E",   x"FC",   x"89",   x"1B", 
  x"79",   x"EB",   x"9E",   x"0C",   x"74",   x"E6",   x"93",   x"01", 
  x"57",   x"C5",   x"B0",   x"22",   x"5A",   x"C8",   x"BD",   x"2F", 
  x"4D",   x"DF",   x"AA",   x"38",   x"40",   x"D2",   x"A7",   x"35", 
  x"0B",   x"99",   x"EC",   x"7E",   x"06",   x"94",   x"E1",   x"73", 
  x"11",   x"83",   x"F6",   x"64",   x"1C",   x"8E",   x"FB",   x"69", 
  x"3F",   x"AD",   x"D8",   x"4A",   x"32",   x"A0",   x"D5",   x"47", 
  x"25",   x"B7",   x"C2",   x"50",   x"28",   x"BA",   x"CF",   x"5D", 
  x"B3",   x"21",   x"54",   x"C6",   x"BE",   x"2C",   x"59",   x"CB", 
  x"A9",   x"3B",   x"4E",   x"DC",   x"A4",   x"36",   x"43",   x"D1", 
  x"87",   x"15",   x"60",   x"F2",   x"8A",   x"18",   x"6D",   x"FF", 
  x"9D",   x"0F",   x"7A",   x"E8",   x"90",   x"02",   x"77",   x"E5", 
  x"DB",   x"49",   x"3C",   x"AE",   x"D6",   x"44",   x"31",   x"A3", 
  x"C1",   x"53",   x"26",   x"B4",   x"CC",   x"5E",   x"2B",   x"B9", 
  x"EF",   x"7D",   x"08",   x"9A",   x"E2",   x"70",   x"05",   x"97", 
  x"F5",   x"67",   x"12",   x"80",   x"F8",   x"6A",   x"1F",   x"8D", 
  x"00",   x"93",   x"E5",   x"76",   x"09",   x"9A",   x"EC",   x"7F", 
  x"12",   x"81",   x"F7",   x"64",   x"1B",   x"88",   x"FE",   x"6D", 
  x"24",   x"B7",   x"C1",   x"52",   x"2D",   x"BE",   x"C8",   x"5B", 
  x"36",   x"A5",   x"D3",   x"40",   x"3F",   x"AC",   x"DA",   x"49", 
  x"48",   x"DB",   x"AD",   x"3E",   x"41",   x"D2",   x"A4",   x"37", 
  x"5A",   x"C9",   x"BF",   x"2C",   x"53",   x"C0",   x"B6",   x"25", 
  x"6C",   x"FF",   x"89",   x"1A",   x"65",   x"F6",   x"80",   x"13", 
  x"7E",   x"ED",   x"9B",   x"08",   x"77",   x"E4",   x"92",   x"01", 
  x"90",   x"03",   x"75",   x"E6",   x"99",   x"0A",   x"7C",   x"EF", 
  x"82",   x"11",   x"67",   x"F4",   x"8B",   x"18",   x"6E",   x"FD", 
  x"B4",   x"27",   x"51",   x"C2",   x"BD",   x"2E",   x"58",   x"CB", 
  x"A6",   x"35",   x"43",   x"D0",   x"AF",   x"3C",   x"4A",   x"D9", 
  x"D8",   x"4B",   x"3D",   x"AE",   x"D1",   x"42",   x"34",   x"A7", 
  x"CA",   x"59",   x"2F",   x"BC",   x"C3",   x"50",   x"26",   x"B5", 
  x"FC",   x"6F",   x"19",   x"8A",   x"F5",   x"66",   x"10",   x"83", 
  x"EE",   x"7D",   x"0B",   x"98",   x"E7",   x"74",   x"02",   x"91", 
  x"E3",   x"70",   x"06",   x"95",   x"EA",   x"79",   x"0F",   x"9C", 
  x"F1",   x"62",   x"14",   x"87",   x"F8",   x"6B",   x"1D",   x"8E", 
  x"C7",   x"54",   x"22",   x"B1",   x"CE",   x"5D",   x"2B",   x"B8", 
  x"D5",   x"46",   x"30",   x"A3",   x"DC",   x"4F",   x"39",   x"AA", 
  x"AB",   x"38",   x"4E",   x"DD",   x"A2",   x"31",   x"47",   x"D4", 
  x"B9",   x"2A",   x"5C",   x"CF",   x"B0",   x"23",   x"55",   x"C6", 
  x"8F",   x"1C",   x"6A",   x"F9",   x"86",   x"15",   x"63",   x"F0", 
  x"9D",   x"0E",   x"78",   x"EB",   x"94",   x"07",   x"71",   x"E2", 
  x"73",   x"E0",   x"96",   x"05",   x"7A",   x"E9",   x"9F",   x"0C", 
  x"61",   x"F2",   x"84",   x"17",   x"68",   x"FB",   x"8D",   x"1E", 
  x"57",   x"C4",   x"B2",   x"21",   x"5E",   x"CD",   x"BB",   x"28", 
  x"45",   x"D6",   x"A0",   x"33",   x"4C",   x"DF",   x"A9",   x"3A", 
  x"3B",   x"A8",   x"DE",   x"4D",   x"32",   x"A1",   x"D7",   x"44", 
  x"29",   x"BA",   x"CC",   x"5F",   x"20",   x"B3",   x"C5",   x"56", 
  x"1F",   x"8C",   x"FA",   x"69",   x"16",   x"85",   x"F3",   x"60", 
  x"0D",   x"9E",   x"E8",   x"7B",   x"04",   x"97",   x"E1",   x"72", 
  x"00",   x"94",   x"EB",   x"7F",   x"15",   x"81",   x"FE",   x"6A", 
  x"2A",   x"BE",   x"C1",   x"55",   x"3F",   x"AB",   x"D4",   x"40", 
  x"54",   x"C0",   x"BF",   x"2B",   x"41",   x"D5",   x"AA",   x"3E", 
  x"7E",   x"EA",   x"95",   x"01",   x"6B",   x"FF",   x"80",   x"14", 
  x"A8",   x"3C",   x"43",   x"D7",   x"BD",   x"29",   x"56",   x"C2", 
  x"82",   x"16",   x"69",   x"FD",   x"97",   x"03",   x"7C",   x"E8", 
  x"FC",   x"68",   x"17",   x"83",   x"E9",   x"7D",   x"02",   x"96", 
  x"D6",   x"42",   x"3D",   x"A9",   x"C3",   x"57",   x"28",   x"BC", 
  x"93",   x"07",   x"78",   x"EC",   x"86",   x"12",   x"6D",   x"F9", 
  x"B9",   x"2D",   x"52",   x"C6",   x"AC",   x"38",   x"47",   x"D3", 
  x"C7",   x"53",   x"2C",   x"B8",   x"D2",   x"46",   x"39",   x"AD", 
  x"ED",   x"79",   x"06",   x"92",   x"F8",   x"6C",   x"13",   x"87", 
  x"3B",   x"AF",   x"D0",   x"44",   x"2E",   x"BA",   x"C5",   x"51", 
  x"11",   x"85",   x"FA",   x"6E",   x"04",   x"90",   x"EF",   x"7B", 
  x"6F",   x"FB",   x"84",   x"10",   x"7A",   x"EE",   x"91",   x"05", 
  x"45",   x"D1",   x"AE",   x"3A",   x"50",   x"C4",   x"BB",   x"2F", 
  x"E5",   x"71",   x"0E",   x"9A",   x"F0",   x"64",   x"1B",   x"8F", 
  x"CF",   x"5B",   x"24",   x"B0",   x"DA",   x"4E",   x"31",   x"A5", 
  x"B1",   x"25",   x"5A",   x"CE",   x"A4",   x"30",   x"4F",   x"DB", 
  x"9B",   x"0F",   x"70",   x"E4",   x"8E",   x"1A",   x"65",   x"F1", 
  x"4D",   x"D9",   x"A6",   x"32",   x"58",   x"CC",   x"B3",   x"27", 
  x"67",   x"F3",   x"8C",   x"18",   x"72",   x"E6",   x"99",   x"0D", 
  x"19",   x"8D",   x"F2",   x"66",   x"0C",   x"98",   x"E7",   x"73", 
  x"33",   x"A7",   x"D8",   x"4C",   x"26",   x"B2",   x"CD",   x"59", 
  x"76",   x"E2",   x"9D",   x"09",   x"63",   x"F7",   x"88",   x"1C", 
  x"5C",   x"C8",   x"B7",   x"23",   x"49",   x"DD",   x"A2",   x"36", 
  x"22",   x"B6",   x"C9",   x"5D",   x"37",   x"A3",   x"DC",   x"48", 
  x"08",   x"9C",   x"E3",   x"77",   x"1D",   x"89",   x"F6",   x"62", 
  x"DE",   x"4A",   x"35",   x"A1",   x"CB",   x"5F",   x"20",   x"B4", 
  x"F4",   x"60",   x"1F",   x"8B",   x"E1",   x"75",   x"0A",   x"9E", 
  x"8A",   x"1E",   x"61",   x"F5",   x"9F",   x"0B",   x"74",   x"E0", 
  x"A0",   x"34",   x"4B",   x"DF",   x"B5",   x"21",   x"5E",   x"CA", 
  x"00",   x"95",   x"E9",   x"7C",   x"11",   x"84",   x"F8",   x"6D", 
  x"22",   x"B7",   x"CB",   x"5E",   x"33",   x"A6",   x"DA",   x"4F", 
  x"44",   x"D1",   x"AD",   x"38",   x"55",   x"C0",   x"BC",   x"29", 
  x"66",   x"F3",   x"8F",   x"1A",   x"77",   x"E2",   x"9E",   x"0B", 
  x"88",   x"1D",   x"61",   x"F4",   x"99",   x"0C",   x"70",   x"E5", 
  x"AA",   x"3F",   x"43",   x"D6",   x"BB",   x"2E",   x"52",   x"C7", 
  x"CC",   x"59",   x"25",   x"B0",   x"DD",   x"48",   x"34",   x"A1", 
  x"EE",   x"7B",   x"07",   x"92",   x"FF",   x"6A",   x"16",   x"83", 
  x"D3",   x"46",   x"3A",   x"AF",   x"C2",   x"57",   x"2B",   x"BE", 
  x"F1",   x"64",   x"18",   x"8D",   x"E0",   x"75",   x"09",   x"9C", 
  x"97",   x"02",   x"7E",   x"EB",   x"86",   x"13",   x"6F",   x"FA", 
  x"B5",   x"20",   x"5C",   x"C9",   x"A4",   x"31",   x"4D",   x"D8", 
  x"5B",   x"CE",   x"B2",   x"27",   x"4A",   x"DF",   x"A3",   x"36", 
  x"79",   x"EC",   x"90",   x"05",   x"68",   x"FD",   x"81",   x"14", 
  x"1F",   x"8A",   x"F6",   x"63",   x"0E",   x"9B",   x"E7",   x"72", 
  x"3D",   x"A8",   x"D4",   x"41",   x"2C",   x"B9",   x"C5",   x"50", 
  x"65",   x"F0",   x"8C",   x"19",   x"74",   x"E1",   x"9D",   x"08", 
  x"47",   x"D2",   x"AE",   x"3B",   x"56",   x"C3",   x"BF",   x"2A", 
  x"21",   x"B4",   x"C8",   x"5D",   x"30",   x"A5",   x"D9",   x"4C", 
  x"03",   x"96",   x"EA",   x"7F",   x"12",   x"87",   x"FB",   x"6E", 
  x"ED",   x"78",   x"04",   x"91",   x"FC",   x"69",   x"15",   x"80", 
  x"CF",   x"5A",   x"26",   x"B3",   x"DE",   x"4B",   x"37",   x"A2", 
  x"A9",   x"3C",   x"40",   x"D5",   x"B8",   x"2D",   x"51",   x"C4", 
  x"8B",   x"1E",   x"62",   x"F7",   x"9A",   x"0F",   x"73",   x"E6", 
  x"B6",   x"23",   x"5F",   x"CA",   x"A7",   x"32",   x"4E",   x"DB", 
  x"94",   x"01",   x"7D",   x"E8",   x"85",   x"10",   x"6C",   x"F9", 
  x"F2",   x"67",   x"1B",   x"8E",   x"E3",   x"76",   x"0A",   x"9F", 
  x"D0",   x"45",   x"39",   x"AC",   x"C1",   x"54",   x"28",   x"BD", 
  x"3E",   x"AB",   x"D7",   x"42",   x"2F",   x"BA",   x"C6",   x"53", 
  x"1C",   x"89",   x"F5",   x"60",   x"0D",   x"98",   x"E4",   x"71", 
  x"7A",   x"EF",   x"93",   x"06",   x"6B",   x"FE",   x"82",   x"17", 
  x"58",   x"CD",   x"B1",   x"24",   x"49",   x"DC",   x"A0",   x"35", 
  x"00",   x"96",   x"EF",   x"79",   x"1D",   x"8B",   x"F2",   x"64", 
  x"3A",   x"AC",   x"D5",   x"43",   x"27",   x"B1",   x"C8",   x"5E", 
  x"74",   x"E2",   x"9B",   x"0D",   x"69",   x"FF",   x"86",   x"10", 
  x"4E",   x"D8",   x"A1",   x"37",   x"53",   x"C5",   x"BC",   x"2A", 
  x"E8",   x"7E",   x"07",   x"91",   x"F5",   x"63",   x"1A",   x"8C", 
  x"D2",   x"44",   x"3D",   x"AB",   x"CF",   x"59",   x"20",   x"B6", 
  x"9C",   x"0A",   x"73",   x"E5",   x"81",   x"17",   x"6E",   x"F8", 
  x"A6",   x"30",   x"49",   x"DF",   x"BB",   x"2D",   x"54",   x"C2", 
  x"13",   x"85",   x"FC",   x"6A",   x"0E",   x"98",   x"E1",   x"77", 
  x"29",   x"BF",   x"C6",   x"50",   x"34",   x"A2",   x"DB",   x"4D", 
  x"67",   x"F1",   x"88",   x"1E",   x"7A",   x"EC",   x"95",   x"03", 
  x"5D",   x"CB",   x"B2",   x"24",   x"40",   x"D6",   x"AF",   x"39", 
  x"FB",   x"6D",   x"14",   x"82",   x"E6",   x"70",   x"09",   x"9F", 
  x"C1",   x"57",   x"2E",   x"B8",   x"DC",   x"4A",   x"33",   x"A5", 
  x"8F",   x"19",   x"60",   x"F6",   x"92",   x"04",   x"7D",   x"EB", 
  x"B5",   x"23",   x"5A",   x"CC",   x"A8",   x"3E",   x"47",   x"D1", 
  x"26",   x"B0",   x"C9",   x"5F",   x"3B",   x"AD",   x"D4",   x"42", 
  x"1C",   x"8A",   x"F3",   x"65",   x"01",   x"97",   x"EE",   x"78", 
  x"52",   x"C4",   x"BD",   x"2B",   x"4F",   x"D9",   x"A0",   x"36", 
  x"68",   x"FE",   x"87",   x"11",   x"75",   x"E3",   x"9A",   x"0C", 
  x"CE",   x"58",   x"21",   x"B7",   x"D3",   x"45",   x"3C",   x"AA", 
  x"F4",   x"62",   x"1B",   x"8D",   x"E9",   x"7F",   x"06",   x"90", 
  x"BA",   x"2C",   x"55",   x"C3",   x"A7",   x"31",   x"48",   x"DE", 
  x"80",   x"16",   x"6F",   x"F9",   x"9D",   x"0B",   x"72",   x"E4", 
  x"35",   x"A3",   x"DA",   x"4C",   x"28",   x"BE",   x"C7",   x"51", 
  x"0F",   x"99",   x"E0",   x"76",   x"12",   x"84",   x"FD",   x"6B", 
  x"41",   x"D7",   x"AE",   x"38",   x"5C",   x"CA",   x"B3",   x"25", 
  x"7B",   x"ED",   x"94",   x"02",   x"66",   x"F0",   x"89",   x"1F", 
  x"DD",   x"4B",   x"32",   x"A4",   x"C0",   x"56",   x"2F",   x"B9", 
  x"E7",   x"71",   x"08",   x"9E",   x"FA",   x"6C",   x"15",   x"83", 
  x"A9",   x"3F",   x"46",   x"D0",   x"B4",   x"22",   x"5B",   x"CD", 
  x"93",   x"05",   x"7C",   x"EA",   x"8E",   x"18",   x"61",   x"F7", 
  x"00",   x"97",   x"ED",   x"7A",   x"19",   x"8E",   x"F4",   x"63", 
  x"32",   x"A5",   x"DF",   x"48",   x"2B",   x"BC",   x"C6",   x"51", 
  x"64",   x"F3",   x"89",   x"1E",   x"7D",   x"EA",   x"90",   x"07", 
  x"56",   x"C1",   x"BB",   x"2C",   x"4F",   x"D8",   x"A2",   x"35", 
  x"C8",   x"5F",   x"25",   x"B2",   x"D1",   x"46",   x"3C",   x"AB", 
  x"FA",   x"6D",   x"17",   x"80",   x"E3",   x"74",   x"0E",   x"99", 
  x"AC",   x"3B",   x"41",   x"D6",   x"B5",   x"22",   x"58",   x"CF", 
  x"9E",   x"09",   x"73",   x"E4",   x"87",   x"10",   x"6A",   x"FD", 
  x"53",   x"C4",   x"BE",   x"29",   x"4A",   x"DD",   x"A7",   x"30", 
  x"61",   x"F6",   x"8C",   x"1B",   x"78",   x"EF",   x"95",   x"02", 
  x"37",   x"A0",   x"DA",   x"4D",   x"2E",   x"B9",   x"C3",   x"54", 
  x"05",   x"92",   x"E8",   x"7F",   x"1C",   x"8B",   x"F1",   x"66", 
  x"9B",   x"0C",   x"76",   x"E1",   x"82",   x"15",   x"6F",   x"F8", 
  x"A9",   x"3E",   x"44",   x"D3",   x"B0",   x"27",   x"5D",   x"CA", 
  x"FF",   x"68",   x"12",   x"85",   x"E6",   x"71",   x"0B",   x"9C", 
  x"CD",   x"5A",   x"20",   x"B7",   x"D4",   x"43",   x"39",   x"AE", 
  x"A6",   x"31",   x"4B",   x"DC",   x"BF",   x"28",   x"52",   x"C5", 
  x"94",   x"03",   x"79",   x"EE",   x"8D",   x"1A",   x"60",   x"F7", 
  x"C2",   x"55",   x"2F",   x"B8",   x"DB",   x"4C",   x"36",   x"A1", 
  x"F0",   x"67",   x"1D",   x"8A",   x"E9",   x"7E",   x"04",   x"93", 
  x"6E",   x"F9",   x"83",   x"14",   x"77",   x"E0",   x"9A",   x"0D", 
  x"5C",   x"CB",   x"B1",   x"26",   x"45",   x"D2",   x"A8",   x"3F", 
  x"0A",   x"9D",   x"E7",   x"70",   x"13",   x"84",   x"FE",   x"69", 
  x"38",   x"AF",   x"D5",   x"42",   x"21",   x"B6",   x"CC",   x"5B", 
  x"F5",   x"62",   x"18",   x"8F",   x"EC",   x"7B",   x"01",   x"96", 
  x"C7",   x"50",   x"2A",   x"BD",   x"DE",   x"49",   x"33",   x"A4", 
  x"91",   x"06",   x"7C",   x"EB",   x"88",   x"1F",   x"65",   x"F2", 
  x"A3",   x"34",   x"4E",   x"D9",   x"BA",   x"2D",   x"57",   x"C0", 
  x"3D",   x"AA",   x"D0",   x"47",   x"24",   x"B3",   x"C9",   x"5E", 
  x"0F",   x"98",   x"E2",   x"75",   x"16",   x"81",   x"FB",   x"6C", 
  x"59",   x"CE",   x"B4",   x"23",   x"40",   x"D7",   x"AD",   x"3A", 
  x"6B",   x"FC",   x"86",   x"11",   x"72",   x"E5",   x"9F",   x"08", 
  x"00",   x"98",   x"F3",   x"6B",   x"25",   x"BD",   x"D6",   x"4E", 
  x"4A",   x"D2",   x"B9",   x"21",   x"6F",   x"F7",   x"9C",   x"04", 
  x"94",   x"0C",   x"67",   x"FF",   x"B1",   x"29",   x"42",   x"DA", 
  x"DE",   x"46",   x"2D",   x"B5",   x"FB",   x"63",   x"08",   x"90", 
  x"EB",   x"73",   x"18",   x"80",   x"CE",   x"56",   x"3D",   x"A5", 
  x"A1",   x"39",   x"52",   x"CA",   x"84",   x"1C",   x"77",   x"EF", 
  x"7F",   x"E7",   x"8C",   x"14",   x"5A",   x"C2",   x"A9",   x"31", 
  x"35",   x"AD",   x"C6",   x"5E",   x"10",   x"88",   x"E3",   x"7B", 
  x"15",   x"8D",   x"E6",   x"7E",   x"30",   x"A8",   x"C3",   x"5B", 
  x"5F",   x"C7",   x"AC",   x"34",   x"7A",   x"E2",   x"89",   x"11", 
  x"81",   x"19",   x"72",   x"EA",   x"A4",   x"3C",   x"57",   x"CF", 
  x"CB",   x"53",   x"38",   x"A0",   x"EE",   x"76",   x"1D",   x"85", 
  x"FE",   x"66",   x"0D",   x"95",   x"DB",   x"43",   x"28",   x"B0", 
  x"B4",   x"2C",   x"47",   x"DF",   x"91",   x"09",   x"62",   x"FA", 
  x"6A",   x"F2",   x"99",   x"01",   x"4F",   x"D7",   x"BC",   x"24", 
  x"20",   x"B8",   x"D3",   x"4B",   x"05",   x"9D",   x"F6",   x"6E", 
  x"2A",   x"B2",   x"D9",   x"41",   x"0F",   x"97",   x"FC",   x"64", 
  x"60",   x"F8",   x"93",   x"0B",   x"45",   x"DD",   x"B6",   x"2E", 
  x"BE",   x"26",   x"4D",   x"D5",   x"9B",   x"03",   x"68",   x"F0", 
  x"F4",   x"6C",   x"07",   x"9F",   x"D1",   x"49",   x"22",   x"BA", 
  x"C1",   x"59",   x"32",   x"AA",   x"E4",   x"7C",   x"17",   x"8F", 
  x"8B",   x"13",   x"78",   x"E0",   x"AE",   x"36",   x"5D",   x"C5", 
  x"55",   x"CD",   x"A6",   x"3E",   x"70",   x"E8",   x"83",   x"1B", 
  x"1F",   x"87",   x"EC",   x"74",   x"3A",   x"A2",   x"C9",   x"51", 
  x"3F",   x"A7",   x"CC",   x"54",   x"1A",   x"82",   x"E9",   x"71", 
  x"75",   x"ED",   x"86",   x"1E",   x"50",   x"C8",   x"A3",   x"3B", 
  x"AB",   x"33",   x"58",   x"C0",   x"8E",   x"16",   x"7D",   x"E5", 
  x"E1",   x"79",   x"12",   x"8A",   x"C4",   x"5C",   x"37",   x"AF", 
  x"D4",   x"4C",   x"27",   x"BF",   x"F1",   x"69",   x"02",   x"9A", 
  x"9E",   x"06",   x"6D",   x"F5",   x"BB",   x"23",   x"48",   x"D0", 
  x"40",   x"D8",   x"B3",   x"2B",   x"65",   x"FD",   x"96",   x"0E", 
  x"0A",   x"92",   x"F9",   x"61",   x"2F",   x"B7",   x"DC",   x"44", 
  x"00",   x"99",   x"F1",   x"68",   x"21",   x"B8",   x"D0",   x"49", 
  x"42",   x"DB",   x"B3",   x"2A",   x"63",   x"FA",   x"92",   x"0B", 
  x"84",   x"1D",   x"75",   x"EC",   x"A5",   x"3C",   x"54",   x"CD", 
  x"C6",   x"5F",   x"37",   x"AE",   x"E7",   x"7E",   x"16",   x"8F", 
  x"CB",   x"52",   x"3A",   x"A3",   x"EA",   x"73",   x"1B",   x"82", 
  x"89",   x"10",   x"78",   x"E1",   x"A8",   x"31",   x"59",   x"C0", 
  x"4F",   x"D6",   x"BE",   x"27",   x"6E",   x"F7",   x"9F",   x"06", 
  x"0D",   x"94",   x"FC",   x"65",   x"2C",   x"B5",   x"DD",   x"44", 
  x"55",   x"CC",   x"A4",   x"3D",   x"74",   x"ED",   x"85",   x"1C", 
  x"17",   x"8E",   x"E6",   x"7F",   x"36",   x"AF",   x"C7",   x"5E", 
  x"D1",   x"48",   x"20",   x"B9",   x"F0",   x"69",   x"01",   x"98", 
  x"93",   x"0A",   x"62",   x"FB",   x"B2",   x"2B",   x"43",   x"DA", 
  x"9E",   x"07",   x"6F",   x"F6",   x"BF",   x"26",   x"4E",   x"D7", 
  x"DC",   x"45",   x"2D",   x"B4",   x"FD",   x"64",   x"0C",   x"95", 
  x"1A",   x"83",   x"EB",   x"72",   x"3B",   x"A2",   x"CA",   x"53", 
  x"58",   x"C1",   x"A9",   x"30",   x"79",   x"E0",   x"88",   x"11", 
  x"AA",   x"33",   x"5B",   x"C2",   x"8B",   x"12",   x"7A",   x"E3", 
  x"E8",   x"71",   x"19",   x"80",   x"C9",   x"50",   x"38",   x"A1", 
  x"2E",   x"B7",   x"DF",   x"46",   x"0F",   x"96",   x"FE",   x"67", 
  x"6C",   x"F5",   x"9D",   x"04",   x"4D",   x"D4",   x"BC",   x"25", 
  x"61",   x"F8",   x"90",   x"09",   x"40",   x"D9",   x"B1",   x"28", 
  x"23",   x"BA",   x"D2",   x"4B",   x"02",   x"9B",   x"F3",   x"6A", 
  x"E5",   x"7C",   x"14",   x"8D",   x"C4",   x"5D",   x"35",   x"AC", 
  x"A7",   x"3E",   x"56",   x"CF",   x"86",   x"1F",   x"77",   x"EE", 
  x"FF",   x"66",   x"0E",   x"97",   x"DE",   x"47",   x"2F",   x"B6", 
  x"BD",   x"24",   x"4C",   x"D5",   x"9C",   x"05",   x"6D",   x"F4", 
  x"7B",   x"E2",   x"8A",   x"13",   x"5A",   x"C3",   x"AB",   x"32", 
  x"39",   x"A0",   x"C8",   x"51",   x"18",   x"81",   x"E9",   x"70", 
  x"34",   x"AD",   x"C5",   x"5C",   x"15",   x"8C",   x"E4",   x"7D", 
  x"76",   x"EF",   x"87",   x"1E",   x"57",   x"CE",   x"A6",   x"3F", 
  x"B0",   x"29",   x"41",   x"D8",   x"91",   x"08",   x"60",   x"F9", 
  x"F2",   x"6B",   x"03",   x"9A",   x"D3",   x"4A",   x"22",   x"BB", 
  x"00",   x"9A",   x"F7",   x"6D",   x"2D",   x"B7",   x"DA",   x"40", 
  x"5A",   x"C0",   x"AD",   x"37",   x"77",   x"ED",   x"80",   x"1A", 
  x"B4",   x"2E",   x"43",   x"D9",   x"99",   x"03",   x"6E",   x"F4", 
  x"EE",   x"74",   x"19",   x"83",   x"C3",   x"59",   x"34",   x"AE", 
  x"AB",   x"31",   x"5C",   x"C6",   x"86",   x"1C",   x"71",   x"EB", 
  x"F1",   x"6B",   x"06",   x"9C",   x"DC",   x"46",   x"2B",   x"B1", 
  x"1F",   x"85",   x"E8",   x"72",   x"32",   x"A8",   x"C5",   x"5F", 
  x"45",   x"DF",   x"B2",   x"28",   x"68",   x"F2",   x"9F",   x"05", 
  x"95",   x"0F",   x"62",   x"F8",   x"B8",   x"22",   x"4F",   x"D5", 
  x"CF",   x"55",   x"38",   x"A2",   x"E2",   x"78",   x"15",   x"8F", 
  x"21",   x"BB",   x"D6",   x"4C",   x"0C",   x"96",   x"FB",   x"61", 
  x"7B",   x"E1",   x"8C",   x"16",   x"56",   x"CC",   x"A1",   x"3B", 
  x"3E",   x"A4",   x"C9",   x"53",   x"13",   x"89",   x"E4",   x"7E", 
  x"64",   x"FE",   x"93",   x"09",   x"49",   x"D3",   x"BE",   x"24", 
  x"8A",   x"10",   x"7D",   x"E7",   x"A7",   x"3D",   x"50",   x"CA", 
  x"D0",   x"4A",   x"27",   x"BD",   x"FD",   x"67",   x"0A",   x"90", 
  x"E9",   x"73",   x"1E",   x"84",   x"C4",   x"5E",   x"33",   x"A9", 
  x"B3",   x"29",   x"44",   x"DE",   x"9E",   x"04",   x"69",   x"F3", 
  x"5D",   x"C7",   x"AA",   x"30",   x"70",   x"EA",   x"87",   x"1D", 
  x"07",   x"9D",   x"F0",   x"6A",   x"2A",   x"B0",   x"DD",   x"47", 
  x"42",   x"D8",   x"B5",   x"2F",   x"6F",   x"F5",   x"98",   x"02", 
  x"18",   x"82",   x"EF",   x"75",   x"35",   x"AF",   x"C2",   x"58", 
  x"F6",   x"6C",   x"01",   x"9B",   x"DB",   x"41",   x"2C",   x"B6", 
  x"AC",   x"36",   x"5B",   x"C1",   x"81",   x"1B",   x"76",   x"EC", 
  x"7C",   x"E6",   x"8B",   x"11",   x"51",   x"CB",   x"A6",   x"3C", 
  x"26",   x"BC",   x"D1",   x"4B",   x"0B",   x"91",   x"FC",   x"66", 
  x"C8",   x"52",   x"3F",   x"A5",   x"E5",   x"7F",   x"12",   x"88", 
  x"92",   x"08",   x"65",   x"FF",   x"BF",   x"25",   x"48",   x"D2", 
  x"D7",   x"4D",   x"20",   x"BA",   x"FA",   x"60",   x"0D",   x"97", 
  x"8D",   x"17",   x"7A",   x"E0",   x"A0",   x"3A",   x"57",   x"CD", 
  x"63",   x"F9",   x"94",   x"0E",   x"4E",   x"D4",   x"B9",   x"23", 
  x"39",   x"A3",   x"CE",   x"54",   x"14",   x"8E",   x"E3",   x"79", 
  x"00",   x"9B",   x"F5",   x"6E",   x"29",   x"B2",   x"DC",   x"47", 
  x"52",   x"C9",   x"A7",   x"3C",   x"7B",   x"E0",   x"8E",   x"15", 
  x"A4",   x"3F",   x"51",   x"CA",   x"8D",   x"16",   x"78",   x"E3", 
  x"F6",   x"6D",   x"03",   x"98",   x"DF",   x"44",   x"2A",   x"B1", 
  x"8B",   x"10",   x"7E",   x"E5",   x"A2",   x"39",   x"57",   x"CC", 
  x"D9",   x"42",   x"2C",   x"B7",   x"F0",   x"6B",   x"05",   x"9E", 
  x"2F",   x"B4",   x"DA",   x"41",   x"06",   x"9D",   x"F3",   x"68", 
  x"7D",   x"E6",   x"88",   x"13",   x"54",   x"CF",   x"A1",   x"3A", 
  x"D5",   x"4E",   x"20",   x"BB",   x"FC",   x"67",   x"09",   x"92", 
  x"87",   x"1C",   x"72",   x"E9",   x"AE",   x"35",   x"5B",   x"C0", 
  x"71",   x"EA",   x"84",   x"1F",   x"58",   x"C3",   x"AD",   x"36", 
  x"23",   x"B8",   x"D6",   x"4D",   x"0A",   x"91",   x"FF",   x"64", 
  x"5E",   x"C5",   x"AB",   x"30",   x"77",   x"EC",   x"82",   x"19", 
  x"0C",   x"97",   x"F9",   x"62",   x"25",   x"BE",   x"D0",   x"4B", 
  x"FA",   x"61",   x"0F",   x"94",   x"D3",   x"48",   x"26",   x"BD", 
  x"A8",   x"33",   x"5D",   x"C6",   x"81",   x"1A",   x"74",   x"EF", 
  x"69",   x"F2",   x"9C",   x"07",   x"40",   x"DB",   x"B5",   x"2E", 
  x"3B",   x"A0",   x"CE",   x"55",   x"12",   x"89",   x"E7",   x"7C", 
  x"CD",   x"56",   x"38",   x"A3",   x"E4",   x"7F",   x"11",   x"8A", 
  x"9F",   x"04",   x"6A",   x"F1",   x"B6",   x"2D",   x"43",   x"D8", 
  x"E2",   x"79",   x"17",   x"8C",   x"CB",   x"50",   x"3E",   x"A5", 
  x"B0",   x"2B",   x"45",   x"DE",   x"99",   x"02",   x"6C",   x"F7", 
  x"46",   x"DD",   x"B3",   x"28",   x"6F",   x"F4",   x"9A",   x"01", 
  x"14",   x"8F",   x"E1",   x"7A",   x"3D",   x"A6",   x"C8",   x"53", 
  x"BC",   x"27",   x"49",   x"D2",   x"95",   x"0E",   x"60",   x"FB", 
  x"EE",   x"75",   x"1B",   x"80",   x"C7",   x"5C",   x"32",   x"A9", 
  x"18",   x"83",   x"ED",   x"76",   x"31",   x"AA",   x"C4",   x"5F", 
  x"4A",   x"D1",   x"BF",   x"24",   x"63",   x"F8",   x"96",   x"0D", 
  x"37",   x"AC",   x"C2",   x"59",   x"1E",   x"85",   x"EB",   x"70", 
  x"65",   x"FE",   x"90",   x"0B",   x"4C",   x"D7",   x"B9",   x"22", 
  x"93",   x"08",   x"66",   x"FD",   x"BA",   x"21",   x"4F",   x"D4", 
  x"C1",   x"5A",   x"34",   x"AF",   x"E8",   x"73",   x"1D",   x"86", 
  x"00",   x"9C",   x"FB",   x"67",   x"35",   x"A9",   x"CE",   x"52", 
  x"6A",   x"F6",   x"91",   x"0D",   x"5F",   x"C3",   x"A4",   x"38", 
  x"D4",   x"48",   x"2F",   x"B3",   x"E1",   x"7D",   x"1A",   x"86", 
  x"BE",   x"22",   x"45",   x"D9",   x"8B",   x"17",   x"70",   x"EC", 
  x"6B",   x"F7",   x"90",   x"0C",   x"5E",   x"C2",   x"A5",   x"39", 
  x"01",   x"9D",   x"FA",   x"66",   x"34",   x"A8",   x"CF",   x"53", 
  x"BF",   x"23",   x"44",   x"D8",   x"8A",   x"16",   x"71",   x"ED", 
  x"D5",   x"49",   x"2E",   x"B2",   x"E0",   x"7C",   x"1B",   x"87", 
  x"D6",   x"4A",   x"2D",   x"B1",   x"E3",   x"7F",   x"18",   x"84", 
  x"BC",   x"20",   x"47",   x"DB",   x"89",   x"15",   x"72",   x"EE", 
  x"02",   x"9E",   x"F9",   x"65",   x"37",   x"AB",   x"CC",   x"50", 
  x"68",   x"F4",   x"93",   x"0F",   x"5D",   x"C1",   x"A6",   x"3A", 
  x"BD",   x"21",   x"46",   x"DA",   x"88",   x"14",   x"73",   x"EF", 
  x"D7",   x"4B",   x"2C",   x"B0",   x"E2",   x"7E",   x"19",   x"85", 
  x"69",   x"F5",   x"92",   x"0E",   x"5C",   x"C0",   x"A7",   x"3B", 
  x"03",   x"9F",   x"F8",   x"64",   x"36",   x"AA",   x"CD",   x"51", 
  x"6F",   x"F3",   x"94",   x"08",   x"5A",   x"C6",   x"A1",   x"3D", 
  x"05",   x"99",   x"FE",   x"62",   x"30",   x"AC",   x"CB",   x"57", 
  x"BB",   x"27",   x"40",   x"DC",   x"8E",   x"12",   x"75",   x"E9", 
  x"D1",   x"4D",   x"2A",   x"B6",   x"E4",   x"78",   x"1F",   x"83", 
  x"04",   x"98",   x"FF",   x"63",   x"31",   x"AD",   x"CA",   x"56", 
  x"6E",   x"F2",   x"95",   x"09",   x"5B",   x"C7",   x"A0",   x"3C", 
  x"D0",   x"4C",   x"2B",   x"B7",   x"E5",   x"79",   x"1E",   x"82", 
  x"BA",   x"26",   x"41",   x"DD",   x"8F",   x"13",   x"74",   x"E8", 
  x"B9",   x"25",   x"42",   x"DE",   x"8C",   x"10",   x"77",   x"EB", 
  x"D3",   x"4F",   x"28",   x"B4",   x"E6",   x"7A",   x"1D",   x"81", 
  x"6D",   x"F1",   x"96",   x"0A",   x"58",   x"C4",   x"A3",   x"3F", 
  x"07",   x"9B",   x"FC",   x"60",   x"32",   x"AE",   x"C9",   x"55", 
  x"D2",   x"4E",   x"29",   x"B5",   x"E7",   x"7B",   x"1C",   x"80", 
  x"B8",   x"24",   x"43",   x"DF",   x"8D",   x"11",   x"76",   x"EA", 
  x"06",   x"9A",   x"FD",   x"61",   x"33",   x"AF",   x"C8",   x"54", 
  x"6C",   x"F0",   x"97",   x"0B",   x"59",   x"C5",   x"A2",   x"3E", 
  x"00",   x"9D",   x"F9",   x"64",   x"31",   x"AC",   x"C8",   x"55", 
  x"62",   x"FF",   x"9B",   x"06",   x"53",   x"CE",   x"AA",   x"37", 
  x"C4",   x"59",   x"3D",   x"A0",   x"F5",   x"68",   x"0C",   x"91", 
  x"A6",   x"3B",   x"5F",   x"C2",   x"97",   x"0A",   x"6E",   x"F3", 
  x"4B",   x"D6",   x"B2",   x"2F",   x"7A",   x"E7",   x"83",   x"1E", 
  x"29",   x"B4",   x"D0",   x"4D",   x"18",   x"85",   x"E1",   x"7C", 
  x"8F",   x"12",   x"76",   x"EB",   x"BE",   x"23",   x"47",   x"DA", 
  x"ED",   x"70",   x"14",   x"89",   x"DC",   x"41",   x"25",   x"B8", 
  x"96",   x"0B",   x"6F",   x"F2",   x"A7",   x"3A",   x"5E",   x"C3", 
  x"F4",   x"69",   x"0D",   x"90",   x"C5",   x"58",   x"3C",   x"A1", 
  x"52",   x"CF",   x"AB",   x"36",   x"63",   x"FE",   x"9A",   x"07", 
  x"30",   x"AD",   x"C9",   x"54",   x"01",   x"9C",   x"F8",   x"65", 
  x"DD",   x"40",   x"24",   x"B9",   x"EC",   x"71",   x"15",   x"88", 
  x"BF",   x"22",   x"46",   x"DB",   x"8E",   x"13",   x"77",   x"EA", 
  x"19",   x"84",   x"E0",   x"7D",   x"28",   x"B5",   x"D1",   x"4C", 
  x"7B",   x"E6",   x"82",   x"1F",   x"4A",   x"D7",   x"B3",   x"2E", 
  x"EF",   x"72",   x"16",   x"8B",   x"DE",   x"43",   x"27",   x"BA", 
  x"8D",   x"10",   x"74",   x"E9",   x"BC",   x"21",   x"45",   x"D8", 
  x"2B",   x"B6",   x"D2",   x"4F",   x"1A",   x"87",   x"E3",   x"7E", 
  x"49",   x"D4",   x"B0",   x"2D",   x"78",   x"E5",   x"81",   x"1C", 
  x"A4",   x"39",   x"5D",   x"C0",   x"95",   x"08",   x"6C",   x"F1", 
  x"C6",   x"5B",   x"3F",   x"A2",   x"F7",   x"6A",   x"0E",   x"93", 
  x"60",   x"FD",   x"99",   x"04",   x"51",   x"CC",   x"A8",   x"35", 
  x"02",   x"9F",   x"FB",   x"66",   x"33",   x"AE",   x"CA",   x"57", 
  x"79",   x"E4",   x"80",   x"1D",   x"48",   x"D5",   x"B1",   x"2C", 
  x"1B",   x"86",   x"E2",   x"7F",   x"2A",   x"B7",   x"D3",   x"4E", 
  x"BD",   x"20",   x"44",   x"D9",   x"8C",   x"11",   x"75",   x"E8", 
  x"DF",   x"42",   x"26",   x"BB",   x"EE",   x"73",   x"17",   x"8A", 
  x"32",   x"AF",   x"CB",   x"56",   x"03",   x"9E",   x"FA",   x"67", 
  x"50",   x"CD",   x"A9",   x"34",   x"61",   x"FC",   x"98",   x"05", 
  x"F6",   x"6B",   x"0F",   x"92",   x"C7",   x"5A",   x"3E",   x"A3", 
  x"94",   x"09",   x"6D",   x"F0",   x"A5",   x"38",   x"5C",   x"C1", 
  x"00",   x"9E",   x"FF",   x"61",   x"3D",   x"A3",   x"C2",   x"5C", 
  x"7A",   x"E4",   x"85",   x"1B",   x"47",   x"D9",   x"B8",   x"26", 
  x"F4",   x"6A",   x"0B",   x"95",   x"C9",   x"57",   x"36",   x"A8", 
  x"8E",   x"10",   x"71",   x"EF",   x"B3",   x"2D",   x"4C",   x"D2", 
  x"2B",   x"B5",   x"D4",   x"4A",   x"16",   x"88",   x"E9",   x"77", 
  x"51",   x"CF",   x"AE",   x"30",   x"6C",   x"F2",   x"93",   x"0D", 
  x"DF",   x"41",   x"20",   x"BE",   x"E2",   x"7C",   x"1D",   x"83", 
  x"A5",   x"3B",   x"5A",   x"C4",   x"98",   x"06",   x"67",   x"F9", 
  x"56",   x"C8",   x"A9",   x"37",   x"6B",   x"F5",   x"94",   x"0A", 
  x"2C",   x"B2",   x"D3",   x"4D",   x"11",   x"8F",   x"EE",   x"70", 
  x"A2",   x"3C",   x"5D",   x"C3",   x"9F",   x"01",   x"60",   x"FE", 
  x"D8",   x"46",   x"27",   x"B9",   x"E5",   x"7B",   x"1A",   x"84", 
  x"7D",   x"E3",   x"82",   x"1C",   x"40",   x"DE",   x"BF",   x"21", 
  x"07",   x"99",   x"F8",   x"66",   x"3A",   x"A4",   x"C5",   x"5B", 
  x"89",   x"17",   x"76",   x"E8",   x"B4",   x"2A",   x"4B",   x"D5", 
  x"F3",   x"6D",   x"0C",   x"92",   x"CE",   x"50",   x"31",   x"AF", 
  x"AC",   x"32",   x"53",   x"CD",   x"91",   x"0F",   x"6E",   x"F0", 
  x"D6",   x"48",   x"29",   x"B7",   x"EB",   x"75",   x"14",   x"8A", 
  x"58",   x"C6",   x"A7",   x"39",   x"65",   x"FB",   x"9A",   x"04", 
  x"22",   x"BC",   x"DD",   x"43",   x"1F",   x"81",   x"E0",   x"7E", 
  x"87",   x"19",   x"78",   x"E6",   x"BA",   x"24",   x"45",   x"DB", 
  x"FD",   x"63",   x"02",   x"9C",   x"C0",   x"5E",   x"3F",   x"A1", 
  x"73",   x"ED",   x"8C",   x"12",   x"4E",   x"D0",   x"B1",   x"2F", 
  x"09",   x"97",   x"F6",   x"68",   x"34",   x"AA",   x"CB",   x"55", 
  x"FA",   x"64",   x"05",   x"9B",   x"C7",   x"59",   x"38",   x"A6", 
  x"80",   x"1E",   x"7F",   x"E1",   x"BD",   x"23",   x"42",   x"DC", 
  x"0E",   x"90",   x"F1",   x"6F",   x"33",   x"AD",   x"CC",   x"52", 
  x"74",   x"EA",   x"8B",   x"15",   x"49",   x"D7",   x"B6",   x"28", 
  x"D1",   x"4F",   x"2E",   x"B0",   x"EC",   x"72",   x"13",   x"8D", 
  x"AB",   x"35",   x"54",   x"CA",   x"96",   x"08",   x"69",   x"F7", 
  x"25",   x"BB",   x"DA",   x"44",   x"18",   x"86",   x"E7",   x"79", 
  x"5F",   x"C1",   x"A0",   x"3E",   x"62",   x"FC",   x"9D",   x"03", 
  x"00",   x"9F",   x"FD",   x"62",   x"39",   x"A6",   x"C4",   x"5B", 
  x"72",   x"ED",   x"8F",   x"10",   x"4B",   x"D4",   x"B6",   x"29", 
  x"E4",   x"7B",   x"19",   x"86",   x"DD",   x"42",   x"20",   x"BF", 
  x"96",   x"09",   x"6B",   x"F4",   x"AF",   x"30",   x"52",   x"CD", 
  x"0B",   x"94",   x"F6",   x"69",   x"32",   x"AD",   x"CF",   x"50", 
  x"79",   x"E6",   x"84",   x"1B",   x"40",   x"DF",   x"BD",   x"22", 
  x"EF",   x"70",   x"12",   x"8D",   x"D6",   x"49",   x"2B",   x"B4", 
  x"9D",   x"02",   x"60",   x"FF",   x"A4",   x"3B",   x"59",   x"C6", 
  x"16",   x"89",   x"EB",   x"74",   x"2F",   x"B0",   x"D2",   x"4D", 
  x"64",   x"FB",   x"99",   x"06",   x"5D",   x"C2",   x"A0",   x"3F", 
  x"F2",   x"6D",   x"0F",   x"90",   x"CB",   x"54",   x"36",   x"A9", 
  x"80",   x"1F",   x"7D",   x"E2",   x"B9",   x"26",   x"44",   x"DB", 
  x"1D",   x"82",   x"E0",   x"7F",   x"24",   x"BB",   x"D9",   x"46", 
  x"6F",   x"F0",   x"92",   x"0D",   x"56",   x"C9",   x"AB",   x"34", 
  x"F9",   x"66",   x"04",   x"9B",   x"C0",   x"5F",   x"3D",   x"A2", 
  x"8B",   x"14",   x"76",   x"E9",   x"B2",   x"2D",   x"4F",   x"D0", 
  x"2C",   x"B3",   x"D1",   x"4E",   x"15",   x"8A",   x"E8",   x"77", 
  x"5E",   x"C1",   x"A3",   x"3C",   x"67",   x"F8",   x"9A",   x"05", 
  x"C8",   x"57",   x"35",   x"AA",   x"F1",   x"6E",   x"0C",   x"93", 
  x"BA",   x"25",   x"47",   x"D8",   x"83",   x"1C",   x"7E",   x"E1", 
  x"27",   x"B8",   x"DA",   x"45",   x"1E",   x"81",   x"E3",   x"7C", 
  x"55",   x"CA",   x"A8",   x"37",   x"6C",   x"F3",   x"91",   x"0E", 
  x"C3",   x"5C",   x"3E",   x"A1",   x"FA",   x"65",   x"07",   x"98", 
  x"B1",   x"2E",   x"4C",   x"D3",   x"88",   x"17",   x"75",   x"EA", 
  x"3A",   x"A5",   x"C7",   x"58",   x"03",   x"9C",   x"FE",   x"61", 
  x"48",   x"D7",   x"B5",   x"2A",   x"71",   x"EE",   x"8C",   x"13", 
  x"DE",   x"41",   x"23",   x"BC",   x"E7",   x"78",   x"1A",   x"85", 
  x"AC",   x"33",   x"51",   x"CE",   x"95",   x"0A",   x"68",   x"F7", 
  x"31",   x"AE",   x"CC",   x"53",   x"08",   x"97",   x"F5",   x"6A", 
  x"43",   x"DC",   x"BE",   x"21",   x"7A",   x"E5",   x"87",   x"18", 
  x"D5",   x"4A",   x"28",   x"B7",   x"EC",   x"73",   x"11",   x"8E", 
  x"A7",   x"38",   x"5A",   x"C5",   x"9E",   x"01",   x"63",   x"FC", 
  x"00",   x"A0",   x"83",   x"23",   x"C5",   x"65",   x"46",   x"E6", 
  x"49",   x"E9",   x"CA",   x"6A",   x"8C",   x"2C",   x"0F",   x"AF", 
  x"92",   x"32",   x"11",   x"B1",   x"57",   x"F7",   x"D4",   x"74", 
  x"DB",   x"7B",   x"58",   x"F8",   x"1E",   x"BE",   x"9D",   x"3D", 
  x"E7",   x"47",   x"64",   x"C4",   x"22",   x"82",   x"A1",   x"01", 
  x"AE",   x"0E",   x"2D",   x"8D",   x"6B",   x"CB",   x"E8",   x"48", 
  x"75",   x"D5",   x"F6",   x"56",   x"B0",   x"10",   x"33",   x"93", 
  x"3C",   x"9C",   x"BF",   x"1F",   x"F9",   x"59",   x"7A",   x"DA", 
  x"0D",   x"AD",   x"8E",   x"2E",   x"C8",   x"68",   x"4B",   x"EB", 
  x"44",   x"E4",   x"C7",   x"67",   x"81",   x"21",   x"02",   x"A2", 
  x"9F",   x"3F",   x"1C",   x"BC",   x"5A",   x"FA",   x"D9",   x"79", 
  x"D6",   x"76",   x"55",   x"F5",   x"13",   x"B3",   x"90",   x"30", 
  x"EA",   x"4A",   x"69",   x"C9",   x"2F",   x"8F",   x"AC",   x"0C", 
  x"A3",   x"03",   x"20",   x"80",   x"66",   x"C6",   x"E5",   x"45", 
  x"78",   x"D8",   x"FB",   x"5B",   x"BD",   x"1D",   x"3E",   x"9E", 
  x"31",   x"91",   x"B2",   x"12",   x"F4",   x"54",   x"77",   x"D7", 
  x"1A",   x"BA",   x"99",   x"39",   x"DF",   x"7F",   x"5C",   x"FC", 
  x"53",   x"F3",   x"D0",   x"70",   x"96",   x"36",   x"15",   x"B5", 
  x"88",   x"28",   x"0B",   x"AB",   x"4D",   x"ED",   x"CE",   x"6E", 
  x"C1",   x"61",   x"42",   x"E2",   x"04",   x"A4",   x"87",   x"27", 
  x"FD",   x"5D",   x"7E",   x"DE",   x"38",   x"98",   x"BB",   x"1B", 
  x"B4",   x"14",   x"37",   x"97",   x"71",   x"D1",   x"F2",   x"52", 
  x"6F",   x"CF",   x"EC",   x"4C",   x"AA",   x"0A",   x"29",   x"89", 
  x"26",   x"86",   x"A5",   x"05",   x"E3",   x"43",   x"60",   x"C0", 
  x"17",   x"B7",   x"94",   x"34",   x"D2",   x"72",   x"51",   x"F1", 
  x"5E",   x"FE",   x"DD",   x"7D",   x"9B",   x"3B",   x"18",   x"B8", 
  x"85",   x"25",   x"06",   x"A6",   x"40",   x"E0",   x"C3",   x"63", 
  x"CC",   x"6C",   x"4F",   x"EF",   x"09",   x"A9",   x"8A",   x"2A", 
  x"F0",   x"50",   x"73",   x"D3",   x"35",   x"95",   x"B6",   x"16", 
  x"B9",   x"19",   x"3A",   x"9A",   x"7C",   x"DC",   x"FF",   x"5F", 
  x"62",   x"C2",   x"E1",   x"41",   x"A7",   x"07",   x"24",   x"84", 
  x"2B",   x"8B",   x"A8",   x"08",   x"EE",   x"4E",   x"6D",   x"CD", 
  x"00",   x"A1",   x"81",   x"20",   x"C1",   x"60",   x"40",   x"E1", 
  x"41",   x"E0",   x"C0",   x"61",   x"80",   x"21",   x"01",   x"A0", 
  x"82",   x"23",   x"03",   x"A2",   x"43",   x"E2",   x"C2",   x"63", 
  x"C3",   x"62",   x"42",   x"E3",   x"02",   x"A3",   x"83",   x"22", 
  x"C7",   x"66",   x"46",   x"E7",   x"06",   x"A7",   x"87",   x"26", 
  x"86",   x"27",   x"07",   x"A6",   x"47",   x"E6",   x"C6",   x"67", 
  x"45",   x"E4",   x"C4",   x"65",   x"84",   x"25",   x"05",   x"A4", 
  x"04",   x"A5",   x"85",   x"24",   x"C5",   x"64",   x"44",   x"E5", 
  x"4D",   x"EC",   x"CC",   x"6D",   x"8C",   x"2D",   x"0D",   x"AC", 
  x"0C",   x"AD",   x"8D",   x"2C",   x"CD",   x"6C",   x"4C",   x"ED", 
  x"CF",   x"6E",   x"4E",   x"EF",   x"0E",   x"AF",   x"8F",   x"2E", 
  x"8E",   x"2F",   x"0F",   x"AE",   x"4F",   x"EE",   x"CE",   x"6F", 
  x"8A",   x"2B",   x"0B",   x"AA",   x"4B",   x"EA",   x"CA",   x"6B", 
  x"CB",   x"6A",   x"4A",   x"EB",   x"0A",   x"AB",   x"8B",   x"2A", 
  x"08",   x"A9",   x"89",   x"28",   x"C9",   x"68",   x"48",   x"E9", 
  x"49",   x"E8",   x"C8",   x"69",   x"88",   x"29",   x"09",   x"A8", 
  x"9A",   x"3B",   x"1B",   x"BA",   x"5B",   x"FA",   x"DA",   x"7B", 
  x"DB",   x"7A",   x"5A",   x"FB",   x"1A",   x"BB",   x"9B",   x"3A", 
  x"18",   x"B9",   x"99",   x"38",   x"D9",   x"78",   x"58",   x"F9", 
  x"59",   x"F8",   x"D8",   x"79",   x"98",   x"39",   x"19",   x"B8", 
  x"5D",   x"FC",   x"DC",   x"7D",   x"9C",   x"3D",   x"1D",   x"BC", 
  x"1C",   x"BD",   x"9D",   x"3C",   x"DD",   x"7C",   x"5C",   x"FD", 
  x"DF",   x"7E",   x"5E",   x"FF",   x"1E",   x"BF",   x"9F",   x"3E", 
  x"9E",   x"3F",   x"1F",   x"BE",   x"5F",   x"FE",   x"DE",   x"7F", 
  x"D7",   x"76",   x"56",   x"F7",   x"16",   x"B7",   x"97",   x"36", 
  x"96",   x"37",   x"17",   x"B6",   x"57",   x"F6",   x"D6",   x"77", 
  x"55",   x"F4",   x"D4",   x"75",   x"94",   x"35",   x"15",   x"B4", 
  x"14",   x"B5",   x"95",   x"34",   x"D5",   x"74",   x"54",   x"F5", 
  x"10",   x"B1",   x"91",   x"30",   x"D1",   x"70",   x"50",   x"F1", 
  x"51",   x"F0",   x"D0",   x"71",   x"90",   x"31",   x"11",   x"B0", 
  x"92",   x"33",   x"13",   x"B2",   x"53",   x"F2",   x"D2",   x"73", 
  x"D3",   x"72",   x"52",   x"F3",   x"12",   x"B3",   x"93",   x"32", 
  x"00",   x"A2",   x"87",   x"25",   x"CD",   x"6F",   x"4A",   x"E8", 
  x"59",   x"FB",   x"DE",   x"7C",   x"94",   x"36",   x"13",   x"B1", 
  x"B2",   x"10",   x"35",   x"97",   x"7F",   x"DD",   x"F8",   x"5A", 
  x"EB",   x"49",   x"6C",   x"CE",   x"26",   x"84",   x"A1",   x"03", 
  x"A7",   x"05",   x"20",   x"82",   x"6A",   x"C8",   x"ED",   x"4F", 
  x"FE",   x"5C",   x"79",   x"DB",   x"33",   x"91",   x"B4",   x"16", 
  x"15",   x"B7",   x"92",   x"30",   x"D8",   x"7A",   x"5F",   x"FD", 
  x"4C",   x"EE",   x"CB",   x"69",   x"81",   x"23",   x"06",   x"A4", 
  x"8D",   x"2F",   x"0A",   x"A8",   x"40",   x"E2",   x"C7",   x"65", 
  x"D4",   x"76",   x"53",   x"F1",   x"19",   x"BB",   x"9E",   x"3C", 
  x"3F",   x"9D",   x"B8",   x"1A",   x"F2",   x"50",   x"75",   x"D7", 
  x"66",   x"C4",   x"E1",   x"43",   x"AB",   x"09",   x"2C",   x"8E", 
  x"2A",   x"88",   x"AD",   x"0F",   x"E7",   x"45",   x"60",   x"C2", 
  x"73",   x"D1",   x"F4",   x"56",   x"BE",   x"1C",   x"39",   x"9B", 
  x"98",   x"3A",   x"1F",   x"BD",   x"55",   x"F7",   x"D2",   x"70", 
  x"C1",   x"63",   x"46",   x"E4",   x"0C",   x"AE",   x"8B",   x"29", 
  x"D9",   x"7B",   x"5E",   x"FC",   x"14",   x"B6",   x"93",   x"31", 
  x"80",   x"22",   x"07",   x"A5",   x"4D",   x"EF",   x"CA",   x"68", 
  x"6B",   x"C9",   x"EC",   x"4E",   x"A6",   x"04",   x"21",   x"83", 
  x"32",   x"90",   x"B5",   x"17",   x"FF",   x"5D",   x"78",   x"DA", 
  x"7E",   x"DC",   x"F9",   x"5B",   x"B3",   x"11",   x"34",   x"96", 
  x"27",   x"85",   x"A0",   x"02",   x"EA",   x"48",   x"6D",   x"CF", 
  x"CC",   x"6E",   x"4B",   x"E9",   x"01",   x"A3",   x"86",   x"24", 
  x"95",   x"37",   x"12",   x"B0",   x"58",   x"FA",   x"DF",   x"7D", 
  x"54",   x"F6",   x"D3",   x"71",   x"99",   x"3B",   x"1E",   x"BC", 
  x"0D",   x"AF",   x"8A",   x"28",   x"C0",   x"62",   x"47",   x"E5", 
  x"E6",   x"44",   x"61",   x"C3",   x"2B",   x"89",   x"AC",   x"0E", 
  x"BF",   x"1D",   x"38",   x"9A",   x"72",   x"D0",   x"F5",   x"57", 
  x"F3",   x"51",   x"74",   x"D6",   x"3E",   x"9C",   x"B9",   x"1B", 
  x"AA",   x"08",   x"2D",   x"8F",   x"67",   x"C5",   x"E0",   x"42", 
  x"41",   x"E3",   x"C6",   x"64",   x"8C",   x"2E",   x"0B",   x"A9", 
  x"18",   x"BA",   x"9F",   x"3D",   x"D5",   x"77",   x"52",   x"F0", 
  x"00",   x"A3",   x"85",   x"26",   x"C9",   x"6A",   x"4C",   x"EF", 
  x"51",   x"F2",   x"D4",   x"77",   x"98",   x"3B",   x"1D",   x"BE", 
  x"A2",   x"01",   x"27",   x"84",   x"6B",   x"C8",   x"EE",   x"4D", 
  x"F3",   x"50",   x"76",   x"D5",   x"3A",   x"99",   x"BF",   x"1C", 
  x"87",   x"24",   x"02",   x"A1",   x"4E",   x"ED",   x"CB",   x"68", 
  x"D6",   x"75",   x"53",   x"F0",   x"1F",   x"BC",   x"9A",   x"39", 
  x"25",   x"86",   x"A0",   x"03",   x"EC",   x"4F",   x"69",   x"CA", 
  x"74",   x"D7",   x"F1",   x"52",   x"BD",   x"1E",   x"38",   x"9B", 
  x"CD",   x"6E",   x"48",   x"EB",   x"04",   x"A7",   x"81",   x"22", 
  x"9C",   x"3F",   x"19",   x"BA",   x"55",   x"F6",   x"D0",   x"73", 
  x"6F",   x"CC",   x"EA",   x"49",   x"A6",   x"05",   x"23",   x"80", 
  x"3E",   x"9D",   x"BB",   x"18",   x"F7",   x"54",   x"72",   x"D1", 
  x"4A",   x"E9",   x"CF",   x"6C",   x"83",   x"20",   x"06",   x"A5", 
  x"1B",   x"B8",   x"9E",   x"3D",   x"D2",   x"71",   x"57",   x"F4", 
  x"E8",   x"4B",   x"6D",   x"CE",   x"21",   x"82",   x"A4",   x"07", 
  x"B9",   x"1A",   x"3C",   x"9F",   x"70",   x"D3",   x"F5",   x"56", 
  x"59",   x"FA",   x"DC",   x"7F",   x"90",   x"33",   x"15",   x"B6", 
  x"08",   x"AB",   x"8D",   x"2E",   x"C1",   x"62",   x"44",   x"E7", 
  x"FB",   x"58",   x"7E",   x"DD",   x"32",   x"91",   x"B7",   x"14", 
  x"AA",   x"09",   x"2F",   x"8C",   x"63",   x"C0",   x"E6",   x"45", 
  x"DE",   x"7D",   x"5B",   x"F8",   x"17",   x"B4",   x"92",   x"31", 
  x"8F",   x"2C",   x"0A",   x"A9",   x"46",   x"E5",   x"C3",   x"60", 
  x"7C",   x"DF",   x"F9",   x"5A",   x"B5",   x"16",   x"30",   x"93", 
  x"2D",   x"8E",   x"A8",   x"0B",   x"E4",   x"47",   x"61",   x"C2", 
  x"94",   x"37",   x"11",   x"B2",   x"5D",   x"FE",   x"D8",   x"7B", 
  x"C5",   x"66",   x"40",   x"E3",   x"0C",   x"AF",   x"89",   x"2A", 
  x"36",   x"95",   x"B3",   x"10",   x"FF",   x"5C",   x"7A",   x"D9", 
  x"67",   x"C4",   x"E2",   x"41",   x"AE",   x"0D",   x"2B",   x"88", 
  x"13",   x"B0",   x"96",   x"35",   x"DA",   x"79",   x"5F",   x"FC", 
  x"42",   x"E1",   x"C7",   x"64",   x"8B",   x"28",   x"0E",   x"AD", 
  x"B1",   x"12",   x"34",   x"97",   x"78",   x"DB",   x"FD",   x"5E", 
  x"E0",   x"43",   x"65",   x"C6",   x"29",   x"8A",   x"AC",   x"0F", 
  x"00",   x"A4",   x"8B",   x"2F",   x"D5",   x"71",   x"5E",   x"FA", 
  x"69",   x"CD",   x"E2",   x"46",   x"BC",   x"18",   x"37",   x"93", 
  x"D2",   x"76",   x"59",   x"FD",   x"07",   x"A3",   x"8C",   x"28", 
  x"BB",   x"1F",   x"30",   x"94",   x"6E",   x"CA",   x"E5",   x"41", 
  x"67",   x"C3",   x"EC",   x"48",   x"B2",   x"16",   x"39",   x"9D", 
  x"0E",   x"AA",   x"85",   x"21",   x"DB",   x"7F",   x"50",   x"F4", 
  x"B5",   x"11",   x"3E",   x"9A",   x"60",   x"C4",   x"EB",   x"4F", 
  x"DC",   x"78",   x"57",   x"F3",   x"09",   x"AD",   x"82",   x"26", 
  x"CE",   x"6A",   x"45",   x"E1",   x"1B",   x"BF",   x"90",   x"34", 
  x"A7",   x"03",   x"2C",   x"88",   x"72",   x"D6",   x"F9",   x"5D", 
  x"1C",   x"B8",   x"97",   x"33",   x"C9",   x"6D",   x"42",   x"E6", 
  x"75",   x"D1",   x"FE",   x"5A",   x"A0",   x"04",   x"2B",   x"8F", 
  x"A9",   x"0D",   x"22",   x"86",   x"7C",   x"D8",   x"F7",   x"53", 
  x"C0",   x"64",   x"4B",   x"EF",   x"15",   x"B1",   x"9E",   x"3A", 
  x"7B",   x"DF",   x"F0",   x"54",   x"AE",   x"0A",   x"25",   x"81", 
  x"12",   x"B6",   x"99",   x"3D",   x"C7",   x"63",   x"4C",   x"E8", 
  x"5F",   x"FB",   x"D4",   x"70",   x"8A",   x"2E",   x"01",   x"A5", 
  x"36",   x"92",   x"BD",   x"19",   x"E3",   x"47",   x"68",   x"CC", 
  x"8D",   x"29",   x"06",   x"A2",   x"58",   x"FC",   x"D3",   x"77", 
  x"E4",   x"40",   x"6F",   x"CB",   x"31",   x"95",   x"BA",   x"1E", 
  x"38",   x"9C",   x"B3",   x"17",   x"ED",   x"49",   x"66",   x"C2", 
  x"51",   x"F5",   x"DA",   x"7E",   x"84",   x"20",   x"0F",   x"AB", 
  x"EA",   x"4E",   x"61",   x"C5",   x"3F",   x"9B",   x"B4",   x"10", 
  x"83",   x"27",   x"08",   x"AC",   x"56",   x"F2",   x"DD",   x"79", 
  x"91",   x"35",   x"1A",   x"BE",   x"44",   x"E0",   x"CF",   x"6B", 
  x"F8",   x"5C",   x"73",   x"D7",   x"2D",   x"89",   x"A6",   x"02", 
  x"43",   x"E7",   x"C8",   x"6C",   x"96",   x"32",   x"1D",   x"B9", 
  x"2A",   x"8E",   x"A1",   x"05",   x"FF",   x"5B",   x"74",   x"D0", 
  x"F6",   x"52",   x"7D",   x"D9",   x"23",   x"87",   x"A8",   x"0C", 
  x"9F",   x"3B",   x"14",   x"B0",   x"4A",   x"EE",   x"C1",   x"65", 
  x"24",   x"80",   x"AF",   x"0B",   x"F1",   x"55",   x"7A",   x"DE", 
  x"4D",   x"E9",   x"C6",   x"62",   x"98",   x"3C",   x"13",   x"B7", 
  x"00",   x"A5",   x"89",   x"2C",   x"D1",   x"74",   x"58",   x"FD", 
  x"61",   x"C4",   x"E8",   x"4D",   x"B0",   x"15",   x"39",   x"9C", 
  x"C2",   x"67",   x"4B",   x"EE",   x"13",   x"B6",   x"9A",   x"3F", 
  x"A3",   x"06",   x"2A",   x"8F",   x"72",   x"D7",   x"FB",   x"5E", 
  x"47",   x"E2",   x"CE",   x"6B",   x"96",   x"33",   x"1F",   x"BA", 
  x"26",   x"83",   x"AF",   x"0A",   x"F7",   x"52",   x"7E",   x"DB", 
  x"85",   x"20",   x"0C",   x"A9",   x"54",   x"F1",   x"DD",   x"78", 
  x"E4",   x"41",   x"6D",   x"C8",   x"35",   x"90",   x"BC",   x"19", 
  x"8E",   x"2B",   x"07",   x"A2",   x"5F",   x"FA",   x"D6",   x"73", 
  x"EF",   x"4A",   x"66",   x"C3",   x"3E",   x"9B",   x"B7",   x"12", 
  x"4C",   x"E9",   x"C5",   x"60",   x"9D",   x"38",   x"14",   x"B1", 
  x"2D",   x"88",   x"A4",   x"01",   x"FC",   x"59",   x"75",   x"D0", 
  x"C9",   x"6C",   x"40",   x"E5",   x"18",   x"BD",   x"91",   x"34", 
  x"A8",   x"0D",   x"21",   x"84",   x"79",   x"DC",   x"F0",   x"55", 
  x"0B",   x"AE",   x"82",   x"27",   x"DA",   x"7F",   x"53",   x"F6", 
  x"6A",   x"CF",   x"E3",   x"46",   x"BB",   x"1E",   x"32",   x"97", 
  x"DF",   x"7A",   x"56",   x"F3",   x"0E",   x"AB",   x"87",   x"22", 
  x"BE",   x"1B",   x"37",   x"92",   x"6F",   x"CA",   x"E6",   x"43", 
  x"1D",   x"B8",   x"94",   x"31",   x"CC",   x"69",   x"45",   x"E0", 
  x"7C",   x"D9",   x"F5",   x"50",   x"AD",   x"08",   x"24",   x"81", 
  x"98",   x"3D",   x"11",   x"B4",   x"49",   x"EC",   x"C0",   x"65", 
  x"F9",   x"5C",   x"70",   x"D5",   x"28",   x"8D",   x"A1",   x"04", 
  x"5A",   x"FF",   x"D3",   x"76",   x"8B",   x"2E",   x"02",   x"A7", 
  x"3B",   x"9E",   x"B2",   x"17",   x"EA",   x"4F",   x"63",   x"C6", 
  x"51",   x"F4",   x"D8",   x"7D",   x"80",   x"25",   x"09",   x"AC", 
  x"30",   x"95",   x"B9",   x"1C",   x"E1",   x"44",   x"68",   x"CD", 
  x"93",   x"36",   x"1A",   x"BF",   x"42",   x"E7",   x"CB",   x"6E", 
  x"F2",   x"57",   x"7B",   x"DE",   x"23",   x"86",   x"AA",   x"0F", 
  x"16",   x"B3",   x"9F",   x"3A",   x"C7",   x"62",   x"4E",   x"EB", 
  x"77",   x"D2",   x"FE",   x"5B",   x"A6",   x"03",   x"2F",   x"8A", 
  x"D4",   x"71",   x"5D",   x"F8",   x"05",   x"A0",   x"8C",   x"29", 
  x"B5",   x"10",   x"3C",   x"99",   x"64",   x"C1",   x"ED",   x"48", 
  x"00",   x"A6",   x"8F",   x"29",   x"DD",   x"7B",   x"52",   x"F4", 
  x"79",   x"DF",   x"F6",   x"50",   x"A4",   x"02",   x"2B",   x"8D", 
  x"F2",   x"54",   x"7D",   x"DB",   x"2F",   x"89",   x"A0",   x"06", 
  x"8B",   x"2D",   x"04",   x"A2",   x"56",   x"F0",   x"D9",   x"7F", 
  x"27",   x"81",   x"A8",   x"0E",   x"FA",   x"5C",   x"75",   x"D3", 
  x"5E",   x"F8",   x"D1",   x"77",   x"83",   x"25",   x"0C",   x"AA", 
  x"D5",   x"73",   x"5A",   x"FC",   x"08",   x"AE",   x"87",   x"21", 
  x"AC",   x"0A",   x"23",   x"85",   x"71",   x"D7",   x"FE",   x"58", 
  x"4E",   x"E8",   x"C1",   x"67",   x"93",   x"35",   x"1C",   x"BA", 
  x"37",   x"91",   x"B8",   x"1E",   x"EA",   x"4C",   x"65",   x"C3", 
  x"BC",   x"1A",   x"33",   x"95",   x"61",   x"C7",   x"EE",   x"48", 
  x"C5",   x"63",   x"4A",   x"EC",   x"18",   x"BE",   x"97",   x"31", 
  x"69",   x"CF",   x"E6",   x"40",   x"B4",   x"12",   x"3B",   x"9D", 
  x"10",   x"B6",   x"9F",   x"39",   x"CD",   x"6B",   x"42",   x"E4", 
  x"9B",   x"3D",   x"14",   x"B2",   x"46",   x"E0",   x"C9",   x"6F", 
  x"E2",   x"44",   x"6D",   x"CB",   x"3F",   x"99",   x"B0",   x"16", 
  x"9C",   x"3A",   x"13",   x"B5",   x"41",   x"E7",   x"CE",   x"68", 
  x"E5",   x"43",   x"6A",   x"CC",   x"38",   x"9E",   x"B7",   x"11", 
  x"6E",   x"C8",   x"E1",   x"47",   x"B3",   x"15",   x"3C",   x"9A", 
  x"17",   x"B1",   x"98",   x"3E",   x"CA",   x"6C",   x"45",   x"E3", 
  x"BB",   x"1D",   x"34",   x"92",   x"66",   x"C0",   x"E9",   x"4F", 
  x"C2",   x"64",   x"4D",   x"EB",   x"1F",   x"B9",   x"90",   x"36", 
  x"49",   x"EF",   x"C6",   x"60",   x"94",   x"32",   x"1B",   x"BD", 
  x"30",   x"96",   x"BF",   x"19",   x"ED",   x"4B",   x"62",   x"C4", 
  x"D2",   x"74",   x"5D",   x"FB",   x"0F",   x"A9",   x"80",   x"26", 
  x"AB",   x"0D",   x"24",   x"82",   x"76",   x"D0",   x"F9",   x"5F", 
  x"20",   x"86",   x"AF",   x"09",   x"FD",   x"5B",   x"72",   x"D4", 
  x"59",   x"FF",   x"D6",   x"70",   x"84",   x"22",   x"0B",   x"AD", 
  x"F5",   x"53",   x"7A",   x"DC",   x"28",   x"8E",   x"A7",   x"01", 
  x"8C",   x"2A",   x"03",   x"A5",   x"51",   x"F7",   x"DE",   x"78", 
  x"07",   x"A1",   x"88",   x"2E",   x"DA",   x"7C",   x"55",   x"F3", 
  x"7E",   x"D8",   x"F1",   x"57",   x"A3",   x"05",   x"2C",   x"8A", 
  x"00",   x"A7",   x"8D",   x"2A",   x"D9",   x"7E",   x"54",   x"F3", 
  x"71",   x"D6",   x"FC",   x"5B",   x"A8",   x"0F",   x"25",   x"82", 
  x"E2",   x"45",   x"6F",   x"C8",   x"3B",   x"9C",   x"B6",   x"11", 
  x"93",   x"34",   x"1E",   x"B9",   x"4A",   x"ED",   x"C7",   x"60", 
  x"07",   x"A0",   x"8A",   x"2D",   x"DE",   x"79",   x"53",   x"F4", 
  x"76",   x"D1",   x"FB",   x"5C",   x"AF",   x"08",   x"22",   x"85", 
  x"E5",   x"42",   x"68",   x"CF",   x"3C",   x"9B",   x"B1",   x"16", 
  x"94",   x"33",   x"19",   x"BE",   x"4D",   x"EA",   x"C0",   x"67", 
  x"0E",   x"A9",   x"83",   x"24",   x"D7",   x"70",   x"5A",   x"FD", 
  x"7F",   x"D8",   x"F2",   x"55",   x"A6",   x"01",   x"2B",   x"8C", 
  x"EC",   x"4B",   x"61",   x"C6",   x"35",   x"92",   x"B8",   x"1F", 
  x"9D",   x"3A",   x"10",   x"B7",   x"44",   x"E3",   x"C9",   x"6E", 
  x"09",   x"AE",   x"84",   x"23",   x"D0",   x"77",   x"5D",   x"FA", 
  x"78",   x"DF",   x"F5",   x"52",   x"A1",   x"06",   x"2C",   x"8B", 
  x"EB",   x"4C",   x"66",   x"C1",   x"32",   x"95",   x"BF",   x"18", 
  x"9A",   x"3D",   x"17",   x"B0",   x"43",   x"E4",   x"CE",   x"69", 
  x"1C",   x"BB",   x"91",   x"36",   x"C5",   x"62",   x"48",   x"EF", 
  x"6D",   x"CA",   x"E0",   x"47",   x"B4",   x"13",   x"39",   x"9E", 
  x"FE",   x"59",   x"73",   x"D4",   x"27",   x"80",   x"AA",   x"0D", 
  x"8F",   x"28",   x"02",   x"A5",   x"56",   x"F1",   x"DB",   x"7C", 
  x"1B",   x"BC",   x"96",   x"31",   x"C2",   x"65",   x"4F",   x"E8", 
  x"6A",   x"CD",   x"E7",   x"40",   x"B3",   x"14",   x"3E",   x"99", 
  x"F9",   x"5E",   x"74",   x"D3",   x"20",   x"87",   x"AD",   x"0A", 
  x"88",   x"2F",   x"05",   x"A2",   x"51",   x"F6",   x"DC",   x"7B", 
  x"12",   x"B5",   x"9F",   x"38",   x"CB",   x"6C",   x"46",   x"E1", 
  x"63",   x"C4",   x"EE",   x"49",   x"BA",   x"1D",   x"37",   x"90", 
  x"F0",   x"57",   x"7D",   x"DA",   x"29",   x"8E",   x"A4",   x"03", 
  x"81",   x"26",   x"0C",   x"AB",   x"58",   x"FF",   x"D5",   x"72", 
  x"15",   x"B2",   x"98",   x"3F",   x"CC",   x"6B",   x"41",   x"E6", 
  x"64",   x"C3",   x"E9",   x"4E",   x"BD",   x"1A",   x"30",   x"97", 
  x"F7",   x"50",   x"7A",   x"DD",   x"2E",   x"89",   x"A3",   x"04", 
  x"86",   x"21",   x"0B",   x"AC",   x"5F",   x"F8",   x"D2",   x"75", 
  x"00",   x"A8",   x"93",   x"3B",   x"E5",   x"4D",   x"76",   x"DE", 
  x"09",   x"A1",   x"9A",   x"32",   x"EC",   x"44",   x"7F",   x"D7", 
  x"12",   x"BA",   x"81",   x"29",   x"F7",   x"5F",   x"64",   x"CC", 
  x"1B",   x"B3",   x"88",   x"20",   x"FE",   x"56",   x"6D",   x"C5", 
  x"24",   x"8C",   x"B7",   x"1F",   x"C1",   x"69",   x"52",   x"FA", 
  x"2D",   x"85",   x"BE",   x"16",   x"C8",   x"60",   x"5B",   x"F3", 
  x"36",   x"9E",   x"A5",   x"0D",   x"D3",   x"7B",   x"40",   x"E8", 
  x"3F",   x"97",   x"AC",   x"04",   x"DA",   x"72",   x"49",   x"E1", 
  x"48",   x"E0",   x"DB",   x"73",   x"AD",   x"05",   x"3E",   x"96", 
  x"41",   x"E9",   x"D2",   x"7A",   x"A4",   x"0C",   x"37",   x"9F", 
  x"5A",   x"F2",   x"C9",   x"61",   x"BF",   x"17",   x"2C",   x"84", 
  x"53",   x"FB",   x"C0",   x"68",   x"B6",   x"1E",   x"25",   x"8D", 
  x"6C",   x"C4",   x"FF",   x"57",   x"89",   x"21",   x"1A",   x"B2", 
  x"65",   x"CD",   x"F6",   x"5E",   x"80",   x"28",   x"13",   x"BB", 
  x"7E",   x"D6",   x"ED",   x"45",   x"9B",   x"33",   x"08",   x"A0", 
  x"77",   x"DF",   x"E4",   x"4C",   x"92",   x"3A",   x"01",   x"A9", 
  x"90",   x"38",   x"03",   x"AB",   x"75",   x"DD",   x"E6",   x"4E", 
  x"99",   x"31",   x"0A",   x"A2",   x"7C",   x"D4",   x"EF",   x"47", 
  x"82",   x"2A",   x"11",   x"B9",   x"67",   x"CF",   x"F4",   x"5C", 
  x"8B",   x"23",   x"18",   x"B0",   x"6E",   x"C6",   x"FD",   x"55", 
  x"B4",   x"1C",   x"27",   x"8F",   x"51",   x"F9",   x"C2",   x"6A", 
  x"BD",   x"15",   x"2E",   x"86",   x"58",   x"F0",   x"CB",   x"63", 
  x"A6",   x"0E",   x"35",   x"9D",   x"43",   x"EB",   x"D0",   x"78", 
  x"AF",   x"07",   x"3C",   x"94",   x"4A",   x"E2",   x"D9",   x"71", 
  x"D8",   x"70",   x"4B",   x"E3",   x"3D",   x"95",   x"AE",   x"06", 
  x"D1",   x"79",   x"42",   x"EA",   x"34",   x"9C",   x"A7",   x"0F", 
  x"CA",   x"62",   x"59",   x"F1",   x"2F",   x"87",   x"BC",   x"14", 
  x"C3",   x"6B",   x"50",   x"F8",   x"26",   x"8E",   x"B5",   x"1D", 
  x"FC",   x"54",   x"6F",   x"C7",   x"19",   x"B1",   x"8A",   x"22", 
  x"F5",   x"5D",   x"66",   x"CE",   x"10",   x"B8",   x"83",   x"2B", 
  x"EE",   x"46",   x"7D",   x"D5",   x"0B",   x"A3",   x"98",   x"30", 
  x"E7",   x"4F",   x"74",   x"DC",   x"02",   x"AA",   x"91",   x"39", 
  x"00",   x"A9",   x"91",   x"38",   x"E1",   x"48",   x"70",   x"D9", 
  x"01",   x"A8",   x"90",   x"39",   x"E0",   x"49",   x"71",   x"D8", 
  x"02",   x"AB",   x"93",   x"3A",   x"E3",   x"4A",   x"72",   x"DB", 
  x"03",   x"AA",   x"92",   x"3B",   x"E2",   x"4B",   x"73",   x"DA", 
  x"04",   x"AD",   x"95",   x"3C",   x"E5",   x"4C",   x"74",   x"DD", 
  x"05",   x"AC",   x"94",   x"3D",   x"E4",   x"4D",   x"75",   x"DC", 
  x"06",   x"AF",   x"97",   x"3E",   x"E7",   x"4E",   x"76",   x"DF", 
  x"07",   x"AE",   x"96",   x"3F",   x"E6",   x"4F",   x"77",   x"DE", 
  x"08",   x"A1",   x"99",   x"30",   x"E9",   x"40",   x"78",   x"D1", 
  x"09",   x"A0",   x"98",   x"31",   x"E8",   x"41",   x"79",   x"D0", 
  x"0A",   x"A3",   x"9B",   x"32",   x"EB",   x"42",   x"7A",   x"D3", 
  x"0B",   x"A2",   x"9A",   x"33",   x"EA",   x"43",   x"7B",   x"D2", 
  x"0C",   x"A5",   x"9D",   x"34",   x"ED",   x"44",   x"7C",   x"D5", 
  x"0D",   x"A4",   x"9C",   x"35",   x"EC",   x"45",   x"7D",   x"D4", 
  x"0E",   x"A7",   x"9F",   x"36",   x"EF",   x"46",   x"7E",   x"D7", 
  x"0F",   x"A6",   x"9E",   x"37",   x"EE",   x"47",   x"7F",   x"D6", 
  x"10",   x"B9",   x"81",   x"28",   x"F1",   x"58",   x"60",   x"C9", 
  x"11",   x"B8",   x"80",   x"29",   x"F0",   x"59",   x"61",   x"C8", 
  x"12",   x"BB",   x"83",   x"2A",   x"F3",   x"5A",   x"62",   x"CB", 
  x"13",   x"BA",   x"82",   x"2B",   x"F2",   x"5B",   x"63",   x"CA", 
  x"14",   x"BD",   x"85",   x"2C",   x"F5",   x"5C",   x"64",   x"CD", 
  x"15",   x"BC",   x"84",   x"2D",   x"F4",   x"5D",   x"65",   x"CC", 
  x"16",   x"BF",   x"87",   x"2E",   x"F7",   x"5E",   x"66",   x"CF", 
  x"17",   x"BE",   x"86",   x"2F",   x"F6",   x"5F",   x"67",   x"CE", 
  x"18",   x"B1",   x"89",   x"20",   x"F9",   x"50",   x"68",   x"C1", 
  x"19",   x"B0",   x"88",   x"21",   x"F8",   x"51",   x"69",   x"C0", 
  x"1A",   x"B3",   x"8B",   x"22",   x"FB",   x"52",   x"6A",   x"C3", 
  x"1B",   x"B2",   x"8A",   x"23",   x"FA",   x"53",   x"6B",   x"C2", 
  x"1C",   x"B5",   x"8D",   x"24",   x"FD",   x"54",   x"6C",   x"C5", 
  x"1D",   x"B4",   x"8C",   x"25",   x"FC",   x"55",   x"6D",   x"C4", 
  x"1E",   x"B7",   x"8F",   x"26",   x"FF",   x"56",   x"6E",   x"C7", 
  x"1F",   x"B6",   x"8E",   x"27",   x"FE",   x"57",   x"6F",   x"C6", 
  x"00",   x"AA",   x"97",   x"3D",   x"ED",   x"47",   x"7A",   x"D0", 
  x"19",   x"B3",   x"8E",   x"24",   x"F4",   x"5E",   x"63",   x"C9", 
  x"32",   x"98",   x"A5",   x"0F",   x"DF",   x"75",   x"48",   x"E2", 
  x"2B",   x"81",   x"BC",   x"16",   x"C6",   x"6C",   x"51",   x"FB", 
  x"64",   x"CE",   x"F3",   x"59",   x"89",   x"23",   x"1E",   x"B4", 
  x"7D",   x"D7",   x"EA",   x"40",   x"90",   x"3A",   x"07",   x"AD", 
  x"56",   x"FC",   x"C1",   x"6B",   x"BB",   x"11",   x"2C",   x"86", 
  x"4F",   x"E5",   x"D8",   x"72",   x"A2",   x"08",   x"35",   x"9F", 
  x"C8",   x"62",   x"5F",   x"F5",   x"25",   x"8F",   x"B2",   x"18", 
  x"D1",   x"7B",   x"46",   x"EC",   x"3C",   x"96",   x"AB",   x"01", 
  x"FA",   x"50",   x"6D",   x"C7",   x"17",   x"BD",   x"80",   x"2A", 
  x"E3",   x"49",   x"74",   x"DE",   x"0E",   x"A4",   x"99",   x"33", 
  x"AC",   x"06",   x"3B",   x"91",   x"41",   x"EB",   x"D6",   x"7C", 
  x"B5",   x"1F",   x"22",   x"88",   x"58",   x"F2",   x"CF",   x"65", 
  x"9E",   x"34",   x"09",   x"A3",   x"73",   x"D9",   x"E4",   x"4E", 
  x"87",   x"2D",   x"10",   x"BA",   x"6A",   x"C0",   x"FD",   x"57", 
  x"53",   x"F9",   x"C4",   x"6E",   x"BE",   x"14",   x"29",   x"83", 
  x"4A",   x"E0",   x"DD",   x"77",   x"A7",   x"0D",   x"30",   x"9A", 
  x"61",   x"CB",   x"F6",   x"5C",   x"8C",   x"26",   x"1B",   x"B1", 
  x"78",   x"D2",   x"EF",   x"45",   x"95",   x"3F",   x"02",   x"A8", 
  x"37",   x"9D",   x"A0",   x"0A",   x"DA",   x"70",   x"4D",   x"E7", 
  x"2E",   x"84",   x"B9",   x"13",   x"C3",   x"69",   x"54",   x"FE", 
  x"05",   x"AF",   x"92",   x"38",   x"E8",   x"42",   x"7F",   x"D5", 
  x"1C",   x"B6",   x"8B",   x"21",   x"F1",   x"5B",   x"66",   x"CC", 
  x"9B",   x"31",   x"0C",   x"A6",   x"76",   x"DC",   x"E1",   x"4B", 
  x"82",   x"28",   x"15",   x"BF",   x"6F",   x"C5",   x"F8",   x"52", 
  x"A9",   x"03",   x"3E",   x"94",   x"44",   x"EE",   x"D3",   x"79", 
  x"B0",   x"1A",   x"27",   x"8D",   x"5D",   x"F7",   x"CA",   x"60", 
  x"FF",   x"55",   x"68",   x"C2",   x"12",   x"B8",   x"85",   x"2F", 
  x"E6",   x"4C",   x"71",   x"DB",   x"0B",   x"A1",   x"9C",   x"36", 
  x"CD",   x"67",   x"5A",   x"F0",   x"20",   x"8A",   x"B7",   x"1D", 
  x"D4",   x"7E",   x"43",   x"E9",   x"39",   x"93",   x"AE",   x"04", 
  x"00",   x"AB",   x"95",   x"3E",   x"E9",   x"42",   x"7C",   x"D7", 
  x"11",   x"BA",   x"84",   x"2F",   x"F8",   x"53",   x"6D",   x"C6", 
  x"22",   x"89",   x"B7",   x"1C",   x"CB",   x"60",   x"5E",   x"F5", 
  x"33",   x"98",   x"A6",   x"0D",   x"DA",   x"71",   x"4F",   x"E4", 
  x"44",   x"EF",   x"D1",   x"7A",   x"AD",   x"06",   x"38",   x"93", 
  x"55",   x"FE",   x"C0",   x"6B",   x"BC",   x"17",   x"29",   x"82", 
  x"66",   x"CD",   x"F3",   x"58",   x"8F",   x"24",   x"1A",   x"B1", 
  x"77",   x"DC",   x"E2",   x"49",   x"9E",   x"35",   x"0B",   x"A0", 
  x"88",   x"23",   x"1D",   x"B6",   x"61",   x"CA",   x"F4",   x"5F", 
  x"99",   x"32",   x"0C",   x"A7",   x"70",   x"DB",   x"E5",   x"4E", 
  x"AA",   x"01",   x"3F",   x"94",   x"43",   x"E8",   x"D6",   x"7D", 
  x"BB",   x"10",   x"2E",   x"85",   x"52",   x"F9",   x"C7",   x"6C", 
  x"CC",   x"67",   x"59",   x"F2",   x"25",   x"8E",   x"B0",   x"1B", 
  x"DD",   x"76",   x"48",   x"E3",   x"34",   x"9F",   x"A1",   x"0A", 
  x"EE",   x"45",   x"7B",   x"D0",   x"07",   x"AC",   x"92",   x"39", 
  x"FF",   x"54",   x"6A",   x"C1",   x"16",   x"BD",   x"83",   x"28", 
  x"D3",   x"78",   x"46",   x"ED",   x"3A",   x"91",   x"AF",   x"04", 
  x"C2",   x"69",   x"57",   x"FC",   x"2B",   x"80",   x"BE",   x"15", 
  x"F1",   x"5A",   x"64",   x"CF",   x"18",   x"B3",   x"8D",   x"26", 
  x"E0",   x"4B",   x"75",   x"DE",   x"09",   x"A2",   x"9C",   x"37", 
  x"97",   x"3C",   x"02",   x"A9",   x"7E",   x"D5",   x"EB",   x"40", 
  x"86",   x"2D",   x"13",   x"B8",   x"6F",   x"C4",   x"FA",   x"51", 
  x"B5",   x"1E",   x"20",   x"8B",   x"5C",   x"F7",   x"C9",   x"62", 
  x"A4",   x"0F",   x"31",   x"9A",   x"4D",   x"E6",   x"D8",   x"73", 
  x"5B",   x"F0",   x"CE",   x"65",   x"B2",   x"19",   x"27",   x"8C", 
  x"4A",   x"E1",   x"DF",   x"74",   x"A3",   x"08",   x"36",   x"9D", 
  x"79",   x"D2",   x"EC",   x"47",   x"90",   x"3B",   x"05",   x"AE", 
  x"68",   x"C3",   x"FD",   x"56",   x"81",   x"2A",   x"14",   x"BF", 
  x"1F",   x"B4",   x"8A",   x"21",   x"F6",   x"5D",   x"63",   x"C8", 
  x"0E",   x"A5",   x"9B",   x"30",   x"E7",   x"4C",   x"72",   x"D9", 
  x"3D",   x"96",   x"A8",   x"03",   x"D4",   x"7F",   x"41",   x"EA", 
  x"2C",   x"87",   x"B9",   x"12",   x"C5",   x"6E",   x"50",   x"FB", 
  x"00",   x"AC",   x"9B",   x"37",   x"F5",   x"59",   x"6E",   x"C2", 
  x"29",   x"85",   x"B2",   x"1E",   x"DC",   x"70",   x"47",   x"EB", 
  x"52",   x"FE",   x"C9",   x"65",   x"A7",   x"0B",   x"3C",   x"90", 
  x"7B",   x"D7",   x"E0",   x"4C",   x"8E",   x"22",   x"15",   x"B9", 
  x"A4",   x"08",   x"3F",   x"93",   x"51",   x"FD",   x"CA",   x"66", 
  x"8D",   x"21",   x"16",   x"BA",   x"78",   x"D4",   x"E3",   x"4F", 
  x"F6",   x"5A",   x"6D",   x"C1",   x"03",   x"AF",   x"98",   x"34", 
  x"DF",   x"73",   x"44",   x"E8",   x"2A",   x"86",   x"B1",   x"1D", 
  x"8B",   x"27",   x"10",   x"BC",   x"7E",   x"D2",   x"E5",   x"49", 
  x"A2",   x"0E",   x"39",   x"95",   x"57",   x"FB",   x"CC",   x"60", 
  x"D9",   x"75",   x"42",   x"EE",   x"2C",   x"80",   x"B7",   x"1B", 
  x"F0",   x"5C",   x"6B",   x"C7",   x"05",   x"A9",   x"9E",   x"32", 
  x"2F",   x"83",   x"B4",   x"18",   x"DA",   x"76",   x"41",   x"ED", 
  x"06",   x"AA",   x"9D",   x"31",   x"F3",   x"5F",   x"68",   x"C4", 
  x"7D",   x"D1",   x"E6",   x"4A",   x"88",   x"24",   x"13",   x"BF", 
  x"54",   x"F8",   x"CF",   x"63",   x"A1",   x"0D",   x"3A",   x"96", 
  x"D5",   x"79",   x"4E",   x"E2",   x"20",   x"8C",   x"BB",   x"17", 
  x"FC",   x"50",   x"67",   x"CB",   x"09",   x"A5",   x"92",   x"3E", 
  x"87",   x"2B",   x"1C",   x"B0",   x"72",   x"DE",   x"E9",   x"45", 
  x"AE",   x"02",   x"35",   x"99",   x"5B",   x"F7",   x"C0",   x"6C", 
  x"71",   x"DD",   x"EA",   x"46",   x"84",   x"28",   x"1F",   x"B3", 
  x"58",   x"F4",   x"C3",   x"6F",   x"AD",   x"01",   x"36",   x"9A", 
  x"23",   x"8F",   x"B8",   x"14",   x"D6",   x"7A",   x"4D",   x"E1", 
  x"0A",   x"A6",   x"91",   x"3D",   x"FF",   x"53",   x"64",   x"C8", 
  x"5E",   x"F2",   x"C5",   x"69",   x"AB",   x"07",   x"30",   x"9C", 
  x"77",   x"DB",   x"EC",   x"40",   x"82",   x"2E",   x"19",   x"B5", 
  x"0C",   x"A0",   x"97",   x"3B",   x"F9",   x"55",   x"62",   x"CE", 
  x"25",   x"89",   x"BE",   x"12",   x"D0",   x"7C",   x"4B",   x"E7", 
  x"FA",   x"56",   x"61",   x"CD",   x"0F",   x"A3",   x"94",   x"38", 
  x"D3",   x"7F",   x"48",   x"E4",   x"26",   x"8A",   x"BD",   x"11", 
  x"A8",   x"04",   x"33",   x"9F",   x"5D",   x"F1",   x"C6",   x"6A", 
  x"81",   x"2D",   x"1A",   x"B6",   x"74",   x"D8",   x"EF",   x"43", 
  x"00",   x"AD",   x"99",   x"34",   x"F1",   x"5C",   x"68",   x"C5", 
  x"21",   x"8C",   x"B8",   x"15",   x"D0",   x"7D",   x"49",   x"E4", 
  x"42",   x"EF",   x"DB",   x"76",   x"B3",   x"1E",   x"2A",   x"87", 
  x"63",   x"CE",   x"FA",   x"57",   x"92",   x"3F",   x"0B",   x"A6", 
  x"84",   x"29",   x"1D",   x"B0",   x"75",   x"D8",   x"EC",   x"41", 
  x"A5",   x"08",   x"3C",   x"91",   x"54",   x"F9",   x"CD",   x"60", 
  x"C6",   x"6B",   x"5F",   x"F2",   x"37",   x"9A",   x"AE",   x"03", 
  x"E7",   x"4A",   x"7E",   x"D3",   x"16",   x"BB",   x"8F",   x"22", 
  x"CB",   x"66",   x"52",   x"FF",   x"3A",   x"97",   x"A3",   x"0E", 
  x"EA",   x"47",   x"73",   x"DE",   x"1B",   x"B6",   x"82",   x"2F", 
  x"89",   x"24",   x"10",   x"BD",   x"78",   x"D5",   x"E1",   x"4C", 
  x"A8",   x"05",   x"31",   x"9C",   x"59",   x"F4",   x"C0",   x"6D", 
  x"4F",   x"E2",   x"D6",   x"7B",   x"BE",   x"13",   x"27",   x"8A", 
  x"6E",   x"C3",   x"F7",   x"5A",   x"9F",   x"32",   x"06",   x"AB", 
  x"0D",   x"A0",   x"94",   x"39",   x"FC",   x"51",   x"65",   x"C8", 
  x"2C",   x"81",   x"B5",   x"18",   x"DD",   x"70",   x"44",   x"E9", 
  x"55",   x"F8",   x"CC",   x"61",   x"A4",   x"09",   x"3D",   x"90", 
  x"74",   x"D9",   x"ED",   x"40",   x"85",   x"28",   x"1C",   x"B1", 
  x"17",   x"BA",   x"8E",   x"23",   x"E6",   x"4B",   x"7F",   x"D2", 
  x"36",   x"9B",   x"AF",   x"02",   x"C7",   x"6A",   x"5E",   x"F3", 
  x"D1",   x"7C",   x"48",   x"E5",   x"20",   x"8D",   x"B9",   x"14", 
  x"F0",   x"5D",   x"69",   x"C4",   x"01",   x"AC",   x"98",   x"35", 
  x"93",   x"3E",   x"0A",   x"A7",   x"62",   x"CF",   x"FB",   x"56", 
  x"B2",   x"1F",   x"2B",   x"86",   x"43",   x"EE",   x"DA",   x"77", 
  x"9E",   x"33",   x"07",   x"AA",   x"6F",   x"C2",   x"F6",   x"5B", 
  x"BF",   x"12",   x"26",   x"8B",   x"4E",   x"E3",   x"D7",   x"7A", 
  x"DC",   x"71",   x"45",   x"E8",   x"2D",   x"80",   x"B4",   x"19", 
  x"FD",   x"50",   x"64",   x"C9",   x"0C",   x"A1",   x"95",   x"38", 
  x"1A",   x"B7",   x"83",   x"2E",   x"EB",   x"46",   x"72",   x"DF", 
  x"3B",   x"96",   x"A2",   x"0F",   x"CA",   x"67",   x"53",   x"FE", 
  x"58",   x"F5",   x"C1",   x"6C",   x"A9",   x"04",   x"30",   x"9D", 
  x"79",   x"D4",   x"E0",   x"4D",   x"88",   x"25",   x"11",   x"BC", 
  x"00",   x"AE",   x"9F",   x"31",   x"FD",   x"53",   x"62",   x"CC", 
  x"39",   x"97",   x"A6",   x"08",   x"C4",   x"6A",   x"5B",   x"F5", 
  x"72",   x"DC",   x"ED",   x"43",   x"8F",   x"21",   x"10",   x"BE", 
  x"4B",   x"E5",   x"D4",   x"7A",   x"B6",   x"18",   x"29",   x"87", 
  x"E4",   x"4A",   x"7B",   x"D5",   x"19",   x"B7",   x"86",   x"28", 
  x"DD",   x"73",   x"42",   x"EC",   x"20",   x"8E",   x"BF",   x"11", 
  x"96",   x"38",   x"09",   x"A7",   x"6B",   x"C5",   x"F4",   x"5A", 
  x"AF",   x"01",   x"30",   x"9E",   x"52",   x"FC",   x"CD",   x"63", 
  x"0B",   x"A5",   x"94",   x"3A",   x"F6",   x"58",   x"69",   x"C7", 
  x"32",   x"9C",   x"AD",   x"03",   x"CF",   x"61",   x"50",   x"FE", 
  x"79",   x"D7",   x"E6",   x"48",   x"84",   x"2A",   x"1B",   x"B5", 
  x"40",   x"EE",   x"DF",   x"71",   x"BD",   x"13",   x"22",   x"8C", 
  x"EF",   x"41",   x"70",   x"DE",   x"12",   x"BC",   x"8D",   x"23", 
  x"D6",   x"78",   x"49",   x"E7",   x"2B",   x"85",   x"B4",   x"1A", 
  x"9D",   x"33",   x"02",   x"AC",   x"60",   x"CE",   x"FF",   x"51", 
  x"A4",   x"0A",   x"3B",   x"95",   x"59",   x"F7",   x"C6",   x"68", 
  x"16",   x"B8",   x"89",   x"27",   x"EB",   x"45",   x"74",   x"DA", 
  x"2F",   x"81",   x"B0",   x"1E",   x"D2",   x"7C",   x"4D",   x"E3", 
  x"64",   x"CA",   x"FB",   x"55",   x"99",   x"37",   x"06",   x"A8", 
  x"5D",   x"F3",   x"C2",   x"6C",   x"A0",   x"0E",   x"3F",   x"91", 
  x"F2",   x"5C",   x"6D",   x"C3",   x"0F",   x"A1",   x"90",   x"3E", 
  x"CB",   x"65",   x"54",   x"FA",   x"36",   x"98",   x"A9",   x"07", 
  x"80",   x"2E",   x"1F",   x"B1",   x"7D",   x"D3",   x"E2",   x"4C", 
  x"B9",   x"17",   x"26",   x"88",   x"44",   x"EA",   x"DB",   x"75", 
  x"1D",   x"B3",   x"82",   x"2C",   x"E0",   x"4E",   x"7F",   x"D1", 
  x"24",   x"8A",   x"BB",   x"15",   x"D9",   x"77",   x"46",   x"E8", 
  x"6F",   x"C1",   x"F0",   x"5E",   x"92",   x"3C",   x"0D",   x"A3", 
  x"56",   x"F8",   x"C9",   x"67",   x"AB",   x"05",   x"34",   x"9A", 
  x"F9",   x"57",   x"66",   x"C8",   x"04",   x"AA",   x"9B",   x"35", 
  x"C0",   x"6E",   x"5F",   x"F1",   x"3D",   x"93",   x"A2",   x"0C", 
  x"8B",   x"25",   x"14",   x"BA",   x"76",   x"D8",   x"E9",   x"47", 
  x"B2",   x"1C",   x"2D",   x"83",   x"4F",   x"E1",   x"D0",   x"7E", 
  x"00",   x"AF",   x"9D",   x"32",   x"F9",   x"56",   x"64",   x"CB", 
  x"31",   x"9E",   x"AC",   x"03",   x"C8",   x"67",   x"55",   x"FA", 
  x"62",   x"CD",   x"FF",   x"50",   x"9B",   x"34",   x"06",   x"A9", 
  x"53",   x"FC",   x"CE",   x"61",   x"AA",   x"05",   x"37",   x"98", 
  x"C4",   x"6B",   x"59",   x"F6",   x"3D",   x"92",   x"A0",   x"0F", 
  x"F5",   x"5A",   x"68",   x"C7",   x"0C",   x"A3",   x"91",   x"3E", 
  x"A6",   x"09",   x"3B",   x"94",   x"5F",   x"F0",   x"C2",   x"6D", 
  x"97",   x"38",   x"0A",   x"A5",   x"6E",   x"C1",   x"F3",   x"5C", 
  x"4B",   x"E4",   x"D6",   x"79",   x"B2",   x"1D",   x"2F",   x"80", 
  x"7A",   x"D5",   x"E7",   x"48",   x"83",   x"2C",   x"1E",   x"B1", 
  x"29",   x"86",   x"B4",   x"1B",   x"D0",   x"7F",   x"4D",   x"E2", 
  x"18",   x"B7",   x"85",   x"2A",   x"E1",   x"4E",   x"7C",   x"D3", 
  x"8F",   x"20",   x"12",   x"BD",   x"76",   x"D9",   x"EB",   x"44", 
  x"BE",   x"11",   x"23",   x"8C",   x"47",   x"E8",   x"DA",   x"75", 
  x"ED",   x"42",   x"70",   x"DF",   x"14",   x"BB",   x"89",   x"26", 
  x"DC",   x"73",   x"41",   x"EE",   x"25",   x"8A",   x"B8",   x"17", 
  x"96",   x"39",   x"0B",   x"A4",   x"6F",   x"C0",   x"F2",   x"5D", 
  x"A7",   x"08",   x"3A",   x"95",   x"5E",   x"F1",   x"C3",   x"6C", 
  x"F4",   x"5B",   x"69",   x"C6",   x"0D",   x"A2",   x"90",   x"3F", 
  x"C5",   x"6A",   x"58",   x"F7",   x"3C",   x"93",   x"A1",   x"0E", 
  x"52",   x"FD",   x"CF",   x"60",   x"AB",   x"04",   x"36",   x"99", 
  x"63",   x"CC",   x"FE",   x"51",   x"9A",   x"35",   x"07",   x"A8", 
  x"30",   x"9F",   x"AD",   x"02",   x"C9",   x"66",   x"54",   x"FB", 
  x"01",   x"AE",   x"9C",   x"33",   x"F8",   x"57",   x"65",   x"CA", 
  x"DD",   x"72",   x"40",   x"EF",   x"24",   x"8B",   x"B9",   x"16", 
  x"EC",   x"43",   x"71",   x"DE",   x"15",   x"BA",   x"88",   x"27", 
  x"BF",   x"10",   x"22",   x"8D",   x"46",   x"E9",   x"DB",   x"74", 
  x"8E",   x"21",   x"13",   x"BC",   x"77",   x"D8",   x"EA",   x"45", 
  x"19",   x"B6",   x"84",   x"2B",   x"E0",   x"4F",   x"7D",   x"D2", 
  x"28",   x"87",   x"B5",   x"1A",   x"D1",   x"7E",   x"4C",   x"E3", 
  x"7B",   x"D4",   x"E6",   x"49",   x"82",   x"2D",   x"1F",   x"B0", 
  x"4A",   x"E5",   x"D7",   x"78",   x"B3",   x"1C",   x"2E",   x"81", 
  x"00",   x"B0",   x"A3",   x"13",   x"85",   x"35",   x"26",   x"96", 
  x"C9",   x"79",   x"6A",   x"DA",   x"4C",   x"FC",   x"EF",   x"5F", 
  x"51",   x"E1",   x"F2",   x"42",   x"D4",   x"64",   x"77",   x"C7", 
  x"98",   x"28",   x"3B",   x"8B",   x"1D",   x"AD",   x"BE",   x"0E", 
  x"A2",   x"12",   x"01",   x"B1",   x"27",   x"97",   x"84",   x"34", 
  x"6B",   x"DB",   x"C8",   x"78",   x"EE",   x"5E",   x"4D",   x"FD", 
  x"F3",   x"43",   x"50",   x"E0",   x"76",   x"C6",   x"D5",   x"65", 
  x"3A",   x"8A",   x"99",   x"29",   x"BF",   x"0F",   x"1C",   x"AC", 
  x"87",   x"37",   x"24",   x"94",   x"02",   x"B2",   x"A1",   x"11", 
  x"4E",   x"FE",   x"ED",   x"5D",   x"CB",   x"7B",   x"68",   x"D8", 
  x"D6",   x"66",   x"75",   x"C5",   x"53",   x"E3",   x"F0",   x"40", 
  x"1F",   x"AF",   x"BC",   x"0C",   x"9A",   x"2A",   x"39",   x"89", 
  x"25",   x"95",   x"86",   x"36",   x"A0",   x"10",   x"03",   x"B3", 
  x"EC",   x"5C",   x"4F",   x"FF",   x"69",   x"D9",   x"CA",   x"7A", 
  x"74",   x"C4",   x"D7",   x"67",   x"F1",   x"41",   x"52",   x"E2", 
  x"BD",   x"0D",   x"1E",   x"AE",   x"38",   x"88",   x"9B",   x"2B", 
  x"CD",   x"7D",   x"6E",   x"DE",   x"48",   x"F8",   x"EB",   x"5B", 
  x"04",   x"B4",   x"A7",   x"17",   x"81",   x"31",   x"22",   x"92", 
  x"9C",   x"2C",   x"3F",   x"8F",   x"19",   x"A9",   x"BA",   x"0A", 
  x"55",   x"E5",   x"F6",   x"46",   x"D0",   x"60",   x"73",   x"C3", 
  x"6F",   x"DF",   x"CC",   x"7C",   x"EA",   x"5A",   x"49",   x"F9", 
  x"A6",   x"16",   x"05",   x"B5",   x"23",   x"93",   x"80",   x"30", 
  x"3E",   x"8E",   x"9D",   x"2D",   x"BB",   x"0B",   x"18",   x"A8", 
  x"F7",   x"47",   x"54",   x"E4",   x"72",   x"C2",   x"D1",   x"61", 
  x"4A",   x"FA",   x"E9",   x"59",   x"CF",   x"7F",   x"6C",   x"DC", 
  x"83",   x"33",   x"20",   x"90",   x"06",   x"B6",   x"A5",   x"15", 
  x"1B",   x"AB",   x"B8",   x"08",   x"9E",   x"2E",   x"3D",   x"8D", 
  x"D2",   x"62",   x"71",   x"C1",   x"57",   x"E7",   x"F4",   x"44", 
  x"E8",   x"58",   x"4B",   x"FB",   x"6D",   x"DD",   x"CE",   x"7E", 
  x"21",   x"91",   x"82",   x"32",   x"A4",   x"14",   x"07",   x"B7", 
  x"B9",   x"09",   x"1A",   x"AA",   x"3C",   x"8C",   x"9F",   x"2F", 
  x"70",   x"C0",   x"D3",   x"63",   x"F5",   x"45",   x"56",   x"E6", 
  x"00",   x"B1",   x"A1",   x"10",   x"81",   x"30",   x"20",   x"91", 
  x"C1",   x"70",   x"60",   x"D1",   x"40",   x"F1",   x"E1",   x"50", 
  x"41",   x"F0",   x"E0",   x"51",   x"C0",   x"71",   x"61",   x"D0", 
  x"80",   x"31",   x"21",   x"90",   x"01",   x"B0",   x"A0",   x"11", 
  x"82",   x"33",   x"23",   x"92",   x"03",   x"B2",   x"A2",   x"13", 
  x"43",   x"F2",   x"E2",   x"53",   x"C2",   x"73",   x"63",   x"D2", 
  x"C3",   x"72",   x"62",   x"D3",   x"42",   x"F3",   x"E3",   x"52", 
  x"02",   x"B3",   x"A3",   x"12",   x"83",   x"32",   x"22",   x"93", 
  x"C7",   x"76",   x"66",   x"D7",   x"46",   x"F7",   x"E7",   x"56", 
  x"06",   x"B7",   x"A7",   x"16",   x"87",   x"36",   x"26",   x"97", 
  x"86",   x"37",   x"27",   x"96",   x"07",   x"B6",   x"A6",   x"17", 
  x"47",   x"F6",   x"E6",   x"57",   x"C6",   x"77",   x"67",   x"D6", 
  x"45",   x"F4",   x"E4",   x"55",   x"C4",   x"75",   x"65",   x"D4", 
  x"84",   x"35",   x"25",   x"94",   x"05",   x"B4",   x"A4",   x"15", 
  x"04",   x"B5",   x"A5",   x"14",   x"85",   x"34",   x"24",   x"95", 
  x"C5",   x"74",   x"64",   x"D5",   x"44",   x"F5",   x"E5",   x"54", 
  x"4D",   x"FC",   x"EC",   x"5D",   x"CC",   x"7D",   x"6D",   x"DC", 
  x"8C",   x"3D",   x"2D",   x"9C",   x"0D",   x"BC",   x"AC",   x"1D", 
  x"0C",   x"BD",   x"AD",   x"1C",   x"8D",   x"3C",   x"2C",   x"9D", 
  x"CD",   x"7C",   x"6C",   x"DD",   x"4C",   x"FD",   x"ED",   x"5C", 
  x"CF",   x"7E",   x"6E",   x"DF",   x"4E",   x"FF",   x"EF",   x"5E", 
  x"0E",   x"BF",   x"AF",   x"1E",   x"8F",   x"3E",   x"2E",   x"9F", 
  x"8E",   x"3F",   x"2F",   x"9E",   x"0F",   x"BE",   x"AE",   x"1F", 
  x"4F",   x"FE",   x"EE",   x"5F",   x"CE",   x"7F",   x"6F",   x"DE", 
  x"8A",   x"3B",   x"2B",   x"9A",   x"0B",   x"BA",   x"AA",   x"1B", 
  x"4B",   x"FA",   x"EA",   x"5B",   x"CA",   x"7B",   x"6B",   x"DA", 
  x"CB",   x"7A",   x"6A",   x"DB",   x"4A",   x"FB",   x"EB",   x"5A", 
  x"0A",   x"BB",   x"AB",   x"1A",   x"8B",   x"3A",   x"2A",   x"9B", 
  x"08",   x"B9",   x"A9",   x"18",   x"89",   x"38",   x"28",   x"99", 
  x"C9",   x"78",   x"68",   x"D9",   x"48",   x"F9",   x"E9",   x"58", 
  x"49",   x"F8",   x"E8",   x"59",   x"C8",   x"79",   x"69",   x"D8", 
  x"88",   x"39",   x"29",   x"98",   x"09",   x"B8",   x"A8",   x"19", 
  x"00",   x"B2",   x"A7",   x"15",   x"8D",   x"3F",   x"2A",   x"98", 
  x"D9",   x"6B",   x"7E",   x"CC",   x"54",   x"E6",   x"F3",   x"41", 
  x"71",   x"C3",   x"D6",   x"64",   x"FC",   x"4E",   x"5B",   x"E9", 
  x"A8",   x"1A",   x"0F",   x"BD",   x"25",   x"97",   x"82",   x"30", 
  x"E2",   x"50",   x"45",   x"F7",   x"6F",   x"DD",   x"C8",   x"7A", 
  x"3B",   x"89",   x"9C",   x"2E",   x"B6",   x"04",   x"11",   x"A3", 
  x"93",   x"21",   x"34",   x"86",   x"1E",   x"AC",   x"B9",   x"0B", 
  x"4A",   x"F8",   x"ED",   x"5F",   x"C7",   x"75",   x"60",   x"D2", 
  x"07",   x"B5",   x"A0",   x"12",   x"8A",   x"38",   x"2D",   x"9F", 
  x"DE",   x"6C",   x"79",   x"CB",   x"53",   x"E1",   x"F4",   x"46", 
  x"76",   x"C4",   x"D1",   x"63",   x"FB",   x"49",   x"5C",   x"EE", 
  x"AF",   x"1D",   x"08",   x"BA",   x"22",   x"90",   x"85",   x"37", 
  x"E5",   x"57",   x"42",   x"F0",   x"68",   x"DA",   x"CF",   x"7D", 
  x"3C",   x"8E",   x"9B",   x"29",   x"B1",   x"03",   x"16",   x"A4", 
  x"94",   x"26",   x"33",   x"81",   x"19",   x"AB",   x"BE",   x"0C", 
  x"4D",   x"FF",   x"EA",   x"58",   x"C0",   x"72",   x"67",   x"D5", 
  x"0E",   x"BC",   x"A9",   x"1B",   x"83",   x"31",   x"24",   x"96", 
  x"D7",   x"65",   x"70",   x"C2",   x"5A",   x"E8",   x"FD",   x"4F", 
  x"7F",   x"CD",   x"D8",   x"6A",   x"F2",   x"40",   x"55",   x"E7", 
  x"A6",   x"14",   x"01",   x"B3",   x"2B",   x"99",   x"8C",   x"3E", 
  x"EC",   x"5E",   x"4B",   x"F9",   x"61",   x"D3",   x"C6",   x"74", 
  x"35",   x"87",   x"92",   x"20",   x"B8",   x"0A",   x"1F",   x"AD", 
  x"9D",   x"2F",   x"3A",   x"88",   x"10",   x"A2",   x"B7",   x"05", 
  x"44",   x"F6",   x"E3",   x"51",   x"C9",   x"7B",   x"6E",   x"DC", 
  x"09",   x"BB",   x"AE",   x"1C",   x"84",   x"36",   x"23",   x"91", 
  x"D0",   x"62",   x"77",   x"C5",   x"5D",   x"EF",   x"FA",   x"48", 
  x"78",   x"CA",   x"DF",   x"6D",   x"F5",   x"47",   x"52",   x"E0", 
  x"A1",   x"13",   x"06",   x"B4",   x"2C",   x"9E",   x"8B",   x"39", 
  x"EB",   x"59",   x"4C",   x"FE",   x"66",   x"D4",   x"C1",   x"73", 
  x"32",   x"80",   x"95",   x"27",   x"BF",   x"0D",   x"18",   x"AA", 
  x"9A",   x"28",   x"3D",   x"8F",   x"17",   x"A5",   x"B0",   x"02", 
  x"43",   x"F1",   x"E4",   x"56",   x"CE",   x"7C",   x"69",   x"DB", 
  x"00",   x"B3",   x"A5",   x"16",   x"89",   x"3A",   x"2C",   x"9F", 
  x"D1",   x"62",   x"74",   x"C7",   x"58",   x"EB",   x"FD",   x"4E", 
  x"61",   x"D2",   x"C4",   x"77",   x"E8",   x"5B",   x"4D",   x"FE", 
  x"B0",   x"03",   x"15",   x"A6",   x"39",   x"8A",   x"9C",   x"2F", 
  x"C2",   x"71",   x"67",   x"D4",   x"4B",   x"F8",   x"EE",   x"5D", 
  x"13",   x"A0",   x"B6",   x"05",   x"9A",   x"29",   x"3F",   x"8C", 
  x"A3",   x"10",   x"06",   x"B5",   x"2A",   x"99",   x"8F",   x"3C", 
  x"72",   x"C1",   x"D7",   x"64",   x"FB",   x"48",   x"5E",   x"ED", 
  x"47",   x"F4",   x"E2",   x"51",   x"CE",   x"7D",   x"6B",   x"D8", 
  x"96",   x"25",   x"33",   x"80",   x"1F",   x"AC",   x"BA",   x"09", 
  x"26",   x"95",   x"83",   x"30",   x"AF",   x"1C",   x"0A",   x"B9", 
  x"F7",   x"44",   x"52",   x"E1",   x"7E",   x"CD",   x"DB",   x"68", 
  x"85",   x"36",   x"20",   x"93",   x"0C",   x"BF",   x"A9",   x"1A", 
  x"54",   x"E7",   x"F1",   x"42",   x"DD",   x"6E",   x"78",   x"CB", 
  x"E4",   x"57",   x"41",   x"F2",   x"6D",   x"DE",   x"C8",   x"7B", 
  x"35",   x"86",   x"90",   x"23",   x"BC",   x"0F",   x"19",   x"AA", 
  x"8E",   x"3D",   x"2B",   x"98",   x"07",   x"B4",   x"A2",   x"11", 
  x"5F",   x"EC",   x"FA",   x"49",   x"D6",   x"65",   x"73",   x"C0", 
  x"EF",   x"5C",   x"4A",   x"F9",   x"66",   x"D5",   x"C3",   x"70", 
  x"3E",   x"8D",   x"9B",   x"28",   x"B7",   x"04",   x"12",   x"A1", 
  x"4C",   x"FF",   x"E9",   x"5A",   x"C5",   x"76",   x"60",   x"D3", 
  x"9D",   x"2E",   x"38",   x"8B",   x"14",   x"A7",   x"B1",   x"02", 
  x"2D",   x"9E",   x"88",   x"3B",   x"A4",   x"17",   x"01",   x"B2", 
  x"FC",   x"4F",   x"59",   x"EA",   x"75",   x"C6",   x"D0",   x"63", 
  x"C9",   x"7A",   x"6C",   x"DF",   x"40",   x"F3",   x"E5",   x"56", 
  x"18",   x"AB",   x"BD",   x"0E",   x"91",   x"22",   x"34",   x"87", 
  x"A8",   x"1B",   x"0D",   x"BE",   x"21",   x"92",   x"84",   x"37", 
  x"79",   x"CA",   x"DC",   x"6F",   x"F0",   x"43",   x"55",   x"E6", 
  x"0B",   x"B8",   x"AE",   x"1D",   x"82",   x"31",   x"27",   x"94", 
  x"DA",   x"69",   x"7F",   x"CC",   x"53",   x"E0",   x"F6",   x"45", 
  x"6A",   x"D9",   x"CF",   x"7C",   x"E3",   x"50",   x"46",   x"F5", 
  x"BB",   x"08",   x"1E",   x"AD",   x"32",   x"81",   x"97",   x"24", 
  x"00",   x"B4",   x"AB",   x"1F",   x"95",   x"21",   x"3E",   x"8A", 
  x"E9",   x"5D",   x"42",   x"F6",   x"7C",   x"C8",   x"D7",   x"63", 
  x"11",   x"A5",   x"BA",   x"0E",   x"84",   x"30",   x"2F",   x"9B", 
  x"F8",   x"4C",   x"53",   x"E7",   x"6D",   x"D9",   x"C6",   x"72", 
  x"22",   x"96",   x"89",   x"3D",   x"B7",   x"03",   x"1C",   x"A8", 
  x"CB",   x"7F",   x"60",   x"D4",   x"5E",   x"EA",   x"F5",   x"41", 
  x"33",   x"87",   x"98",   x"2C",   x"A6",   x"12",   x"0D",   x"B9", 
  x"DA",   x"6E",   x"71",   x"C5",   x"4F",   x"FB",   x"E4",   x"50", 
  x"44",   x"F0",   x"EF",   x"5B",   x"D1",   x"65",   x"7A",   x"CE", 
  x"AD",   x"19",   x"06",   x"B2",   x"38",   x"8C",   x"93",   x"27", 
  x"55",   x"E1",   x"FE",   x"4A",   x"C0",   x"74",   x"6B",   x"DF", 
  x"BC",   x"08",   x"17",   x"A3",   x"29",   x"9D",   x"82",   x"36", 
  x"66",   x"D2",   x"CD",   x"79",   x"F3",   x"47",   x"58",   x"EC", 
  x"8F",   x"3B",   x"24",   x"90",   x"1A",   x"AE",   x"B1",   x"05", 
  x"77",   x"C3",   x"DC",   x"68",   x"E2",   x"56",   x"49",   x"FD", 
  x"9E",   x"2A",   x"35",   x"81",   x"0B",   x"BF",   x"A0",   x"14", 
  x"88",   x"3C",   x"23",   x"97",   x"1D",   x"A9",   x"B6",   x"02", 
  x"61",   x"D5",   x"CA",   x"7E",   x"F4",   x"40",   x"5F",   x"EB", 
  x"99",   x"2D",   x"32",   x"86",   x"0C",   x"B8",   x"A7",   x"13", 
  x"70",   x"C4",   x"DB",   x"6F",   x"E5",   x"51",   x"4E",   x"FA", 
  x"AA",   x"1E",   x"01",   x"B5",   x"3F",   x"8B",   x"94",   x"20", 
  x"43",   x"F7",   x"E8",   x"5C",   x"D6",   x"62",   x"7D",   x"C9", 
  x"BB",   x"0F",   x"10",   x"A4",   x"2E",   x"9A",   x"85",   x"31", 
  x"52",   x"E6",   x"F9",   x"4D",   x"C7",   x"73",   x"6C",   x"D8", 
  x"CC",   x"78",   x"67",   x"D3",   x"59",   x"ED",   x"F2",   x"46", 
  x"25",   x"91",   x"8E",   x"3A",   x"B0",   x"04",   x"1B",   x"AF", 
  x"DD",   x"69",   x"76",   x"C2",   x"48",   x"FC",   x"E3",   x"57", 
  x"34",   x"80",   x"9F",   x"2B",   x"A1",   x"15",   x"0A",   x"BE", 
  x"EE",   x"5A",   x"45",   x"F1",   x"7B",   x"CF",   x"D0",   x"64", 
  x"07",   x"B3",   x"AC",   x"18",   x"92",   x"26",   x"39",   x"8D", 
  x"FF",   x"4B",   x"54",   x"E0",   x"6A",   x"DE",   x"C1",   x"75", 
  x"16",   x"A2",   x"BD",   x"09",   x"83",   x"37",   x"28",   x"9C", 
  x"00",   x"B5",   x"A9",   x"1C",   x"91",   x"24",   x"38",   x"8D", 
  x"E1",   x"54",   x"48",   x"FD",   x"70",   x"C5",   x"D9",   x"6C", 
  x"01",   x"B4",   x"A8",   x"1D",   x"90",   x"25",   x"39",   x"8C", 
  x"E0",   x"55",   x"49",   x"FC",   x"71",   x"C4",   x"D8",   x"6D", 
  x"02",   x"B7",   x"AB",   x"1E",   x"93",   x"26",   x"3A",   x"8F", 
  x"E3",   x"56",   x"4A",   x"FF",   x"72",   x"C7",   x"DB",   x"6E", 
  x"03",   x"B6",   x"AA",   x"1F",   x"92",   x"27",   x"3B",   x"8E", 
  x"E2",   x"57",   x"4B",   x"FE",   x"73",   x"C6",   x"DA",   x"6F", 
  x"04",   x"B1",   x"AD",   x"18",   x"95",   x"20",   x"3C",   x"89", 
  x"E5",   x"50",   x"4C",   x"F9",   x"74",   x"C1",   x"DD",   x"68", 
  x"05",   x"B0",   x"AC",   x"19",   x"94",   x"21",   x"3D",   x"88", 
  x"E4",   x"51",   x"4D",   x"F8",   x"75",   x"C0",   x"DC",   x"69", 
  x"06",   x"B3",   x"AF",   x"1A",   x"97",   x"22",   x"3E",   x"8B", 
  x"E7",   x"52",   x"4E",   x"FB",   x"76",   x"C3",   x"DF",   x"6A", 
  x"07",   x"B2",   x"AE",   x"1B",   x"96",   x"23",   x"3F",   x"8A", 
  x"E6",   x"53",   x"4F",   x"FA",   x"77",   x"C2",   x"DE",   x"6B", 
  x"08",   x"BD",   x"A1",   x"14",   x"99",   x"2C",   x"30",   x"85", 
  x"E9",   x"5C",   x"40",   x"F5",   x"78",   x"CD",   x"D1",   x"64", 
  x"09",   x"BC",   x"A0",   x"15",   x"98",   x"2D",   x"31",   x"84", 
  x"E8",   x"5D",   x"41",   x"F4",   x"79",   x"CC",   x"D0",   x"65", 
  x"0A",   x"BF",   x"A3",   x"16",   x"9B",   x"2E",   x"32",   x"87", 
  x"EB",   x"5E",   x"42",   x"F7",   x"7A",   x"CF",   x"D3",   x"66", 
  x"0B",   x"BE",   x"A2",   x"17",   x"9A",   x"2F",   x"33",   x"86", 
  x"EA",   x"5F",   x"43",   x"F6",   x"7B",   x"CE",   x"D2",   x"67", 
  x"0C",   x"B9",   x"A5",   x"10",   x"9D",   x"28",   x"34",   x"81", 
  x"ED",   x"58",   x"44",   x"F1",   x"7C",   x"C9",   x"D5",   x"60", 
  x"0D",   x"B8",   x"A4",   x"11",   x"9C",   x"29",   x"35",   x"80", 
  x"EC",   x"59",   x"45",   x"F0",   x"7D",   x"C8",   x"D4",   x"61", 
  x"0E",   x"BB",   x"A7",   x"12",   x"9F",   x"2A",   x"36",   x"83", 
  x"EF",   x"5A",   x"46",   x"F3",   x"7E",   x"CB",   x"D7",   x"62", 
  x"0F",   x"BA",   x"A6",   x"13",   x"9E",   x"2B",   x"37",   x"82", 
  x"EE",   x"5B",   x"47",   x"F2",   x"7F",   x"CA",   x"D6",   x"63", 
  x"00",   x"B6",   x"AF",   x"19",   x"9D",   x"2B",   x"32",   x"84", 
  x"F9",   x"4F",   x"56",   x"E0",   x"64",   x"D2",   x"CB",   x"7D", 
  x"31",   x"87",   x"9E",   x"28",   x"AC",   x"1A",   x"03",   x"B5", 
  x"C8",   x"7E",   x"67",   x"D1",   x"55",   x"E3",   x"FA",   x"4C", 
  x"62",   x"D4",   x"CD",   x"7B",   x"FF",   x"49",   x"50",   x"E6", 
  x"9B",   x"2D",   x"34",   x"82",   x"06",   x"B0",   x"A9",   x"1F", 
  x"53",   x"E5",   x"FC",   x"4A",   x"CE",   x"78",   x"61",   x"D7", 
  x"AA",   x"1C",   x"05",   x"B3",   x"37",   x"81",   x"98",   x"2E", 
  x"C4",   x"72",   x"6B",   x"DD",   x"59",   x"EF",   x"F6",   x"40", 
  x"3D",   x"8B",   x"92",   x"24",   x"A0",   x"16",   x"0F",   x"B9", 
  x"F5",   x"43",   x"5A",   x"EC",   x"68",   x"DE",   x"C7",   x"71", 
  x"0C",   x"BA",   x"A3",   x"15",   x"91",   x"27",   x"3E",   x"88", 
  x"A6",   x"10",   x"09",   x"BF",   x"3B",   x"8D",   x"94",   x"22", 
  x"5F",   x"E9",   x"F0",   x"46",   x"C2",   x"74",   x"6D",   x"DB", 
  x"97",   x"21",   x"38",   x"8E",   x"0A",   x"BC",   x"A5",   x"13", 
  x"6E",   x"D8",   x"C1",   x"77",   x"F3",   x"45",   x"5C",   x"EA", 
  x"4B",   x"FD",   x"E4",   x"52",   x"D6",   x"60",   x"79",   x"CF", 
  x"B2",   x"04",   x"1D",   x"AB",   x"2F",   x"99",   x"80",   x"36", 
  x"7A",   x"CC",   x"D5",   x"63",   x"E7",   x"51",   x"48",   x"FE", 
  x"83",   x"35",   x"2C",   x"9A",   x"1E",   x"A8",   x"B1",   x"07", 
  x"29",   x"9F",   x"86",   x"30",   x"B4",   x"02",   x"1B",   x"AD", 
  x"D0",   x"66",   x"7F",   x"C9",   x"4D",   x"FB",   x"E2",   x"54", 
  x"18",   x"AE",   x"B7",   x"01",   x"85",   x"33",   x"2A",   x"9C", 
  x"E1",   x"57",   x"4E",   x"F8",   x"7C",   x"CA",   x"D3",   x"65", 
  x"8F",   x"39",   x"20",   x"96",   x"12",   x"A4",   x"BD",   x"0B", 
  x"76",   x"C0",   x"D9",   x"6F",   x"EB",   x"5D",   x"44",   x"F2", 
  x"BE",   x"08",   x"11",   x"A7",   x"23",   x"95",   x"8C",   x"3A", 
  x"47",   x"F1",   x"E8",   x"5E",   x"DA",   x"6C",   x"75",   x"C3", 
  x"ED",   x"5B",   x"42",   x"F4",   x"70",   x"C6",   x"DF",   x"69", 
  x"14",   x"A2",   x"BB",   x"0D",   x"89",   x"3F",   x"26",   x"90", 
  x"DC",   x"6A",   x"73",   x"C5",   x"41",   x"F7",   x"EE",   x"58", 
  x"25",   x"93",   x"8A",   x"3C",   x"B8",   x"0E",   x"17",   x"A1", 
  x"00",   x"B7",   x"AD",   x"1A",   x"99",   x"2E",   x"34",   x"83", 
  x"F1",   x"46",   x"5C",   x"EB",   x"68",   x"DF",   x"C5",   x"72", 
  x"21",   x"96",   x"8C",   x"3B",   x"B8",   x"0F",   x"15",   x"A2", 
  x"D0",   x"67",   x"7D",   x"CA",   x"49",   x"FE",   x"E4",   x"53", 
  x"42",   x"F5",   x"EF",   x"58",   x"DB",   x"6C",   x"76",   x"C1", 
  x"B3",   x"04",   x"1E",   x"A9",   x"2A",   x"9D",   x"87",   x"30", 
  x"63",   x"D4",   x"CE",   x"79",   x"FA",   x"4D",   x"57",   x"E0", 
  x"92",   x"25",   x"3F",   x"88",   x"0B",   x"BC",   x"A6",   x"11", 
  x"84",   x"33",   x"29",   x"9E",   x"1D",   x"AA",   x"B0",   x"07", 
  x"75",   x"C2",   x"D8",   x"6F",   x"EC",   x"5B",   x"41",   x"F6", 
  x"A5",   x"12",   x"08",   x"BF",   x"3C",   x"8B",   x"91",   x"26", 
  x"54",   x"E3",   x"F9",   x"4E",   x"CD",   x"7A",   x"60",   x"D7", 
  x"C6",   x"71",   x"6B",   x"DC",   x"5F",   x"E8",   x"F2",   x"45", 
  x"37",   x"80",   x"9A",   x"2D",   x"AE",   x"19",   x"03",   x"B4", 
  x"E7",   x"50",   x"4A",   x"FD",   x"7E",   x"C9",   x"D3",   x"64", 
  x"16",   x"A1",   x"BB",   x"0C",   x"8F",   x"38",   x"22",   x"95", 
  x"CB",   x"7C",   x"66",   x"D1",   x"52",   x"E5",   x"FF",   x"48", 
  x"3A",   x"8D",   x"97",   x"20",   x"A3",   x"14",   x"0E",   x"B9", 
  x"EA",   x"5D",   x"47",   x"F0",   x"73",   x"C4",   x"DE",   x"69", 
  x"1B",   x"AC",   x"B6",   x"01",   x"82",   x"35",   x"2F",   x"98", 
  x"89",   x"3E",   x"24",   x"93",   x"10",   x"A7",   x"BD",   x"0A", 
  x"78",   x"CF",   x"D5",   x"62",   x"E1",   x"56",   x"4C",   x"FB", 
  x"A8",   x"1F",   x"05",   x"B2",   x"31",   x"86",   x"9C",   x"2B", 
  x"59",   x"EE",   x"F4",   x"43",   x"C0",   x"77",   x"6D",   x"DA", 
  x"4F",   x"F8",   x"E2",   x"55",   x"D6",   x"61",   x"7B",   x"CC", 
  x"BE",   x"09",   x"13",   x"A4",   x"27",   x"90",   x"8A",   x"3D", 
  x"6E",   x"D9",   x"C3",   x"74",   x"F7",   x"40",   x"5A",   x"ED", 
  x"9F",   x"28",   x"32",   x"85",   x"06",   x"B1",   x"AB",   x"1C", 
  x"0D",   x"BA",   x"A0",   x"17",   x"94",   x"23",   x"39",   x"8E", 
  x"FC",   x"4B",   x"51",   x"E6",   x"65",   x"D2",   x"C8",   x"7F", 
  x"2C",   x"9B",   x"81",   x"36",   x"B5",   x"02",   x"18",   x"AF", 
  x"DD",   x"6A",   x"70",   x"C7",   x"44",   x"F3",   x"E9",   x"5E", 
  x"00",   x"B8",   x"B3",   x"0B",   x"A5",   x"1D",   x"16",   x"AE", 
  x"89",   x"31",   x"3A",   x"82",   x"2C",   x"94",   x"9F",   x"27", 
  x"D1",   x"69",   x"62",   x"DA",   x"74",   x"CC",   x"C7",   x"7F", 
  x"58",   x"E0",   x"EB",   x"53",   x"FD",   x"45",   x"4E",   x"F6", 
  x"61",   x"D9",   x"D2",   x"6A",   x"C4",   x"7C",   x"77",   x"CF", 
  x"E8",   x"50",   x"5B",   x"E3",   x"4D",   x"F5",   x"FE",   x"46", 
  x"B0",   x"08",   x"03",   x"BB",   x"15",   x"AD",   x"A6",   x"1E", 
  x"39",   x"81",   x"8A",   x"32",   x"9C",   x"24",   x"2F",   x"97", 
  x"C2",   x"7A",   x"71",   x"C9",   x"67",   x"DF",   x"D4",   x"6C", 
  x"4B",   x"F3",   x"F8",   x"40",   x"EE",   x"56",   x"5D",   x"E5", 
  x"13",   x"AB",   x"A0",   x"18",   x"B6",   x"0E",   x"05",   x"BD", 
  x"9A",   x"22",   x"29",   x"91",   x"3F",   x"87",   x"8C",   x"34", 
  x"A3",   x"1B",   x"10",   x"A8",   x"06",   x"BE",   x"B5",   x"0D", 
  x"2A",   x"92",   x"99",   x"21",   x"8F",   x"37",   x"3C",   x"84", 
  x"72",   x"CA",   x"C1",   x"79",   x"D7",   x"6F",   x"64",   x"DC", 
  x"FB",   x"43",   x"48",   x"F0",   x"5E",   x"E6",   x"ED",   x"55", 
  x"47",   x"FF",   x"F4",   x"4C",   x"E2",   x"5A",   x"51",   x"E9", 
  x"CE",   x"76",   x"7D",   x"C5",   x"6B",   x"D3",   x"D8",   x"60", 
  x"96",   x"2E",   x"25",   x"9D",   x"33",   x"8B",   x"80",   x"38", 
  x"1F",   x"A7",   x"AC",   x"14",   x"BA",   x"02",   x"09",   x"B1", 
  x"26",   x"9E",   x"95",   x"2D",   x"83",   x"3B",   x"30",   x"88", 
  x"AF",   x"17",   x"1C",   x"A4",   x"0A",   x"B2",   x"B9",   x"01", 
  x"F7",   x"4F",   x"44",   x"FC",   x"52",   x"EA",   x"E1",   x"59", 
  x"7E",   x"C6",   x"CD",   x"75",   x"DB",   x"63",   x"68",   x"D0", 
  x"85",   x"3D",   x"36",   x"8E",   x"20",   x"98",   x"93",   x"2B", 
  x"0C",   x"B4",   x"BF",   x"07",   x"A9",   x"11",   x"1A",   x"A2", 
  x"54",   x"EC",   x"E7",   x"5F",   x"F1",   x"49",   x"42",   x"FA", 
  x"DD",   x"65",   x"6E",   x"D6",   x"78",   x"C0",   x"CB",   x"73", 
  x"E4",   x"5C",   x"57",   x"EF",   x"41",   x"F9",   x"F2",   x"4A", 
  x"6D",   x"D5",   x"DE",   x"66",   x"C8",   x"70",   x"7B",   x"C3", 
  x"35",   x"8D",   x"86",   x"3E",   x"90",   x"28",   x"23",   x"9B", 
  x"BC",   x"04",   x"0F",   x"B7",   x"19",   x"A1",   x"AA",   x"12", 
  x"00",   x"B9",   x"B1",   x"08",   x"A1",   x"18",   x"10",   x"A9", 
  x"81",   x"38",   x"30",   x"89",   x"20",   x"99",   x"91",   x"28", 
  x"C1",   x"78",   x"70",   x"C9",   x"60",   x"D9",   x"D1",   x"68", 
  x"40",   x"F9",   x"F1",   x"48",   x"E1",   x"58",   x"50",   x"E9", 
  x"41",   x"F8",   x"F0",   x"49",   x"E0",   x"59",   x"51",   x"E8", 
  x"C0",   x"79",   x"71",   x"C8",   x"61",   x"D8",   x"D0",   x"69", 
  x"80",   x"39",   x"31",   x"88",   x"21",   x"98",   x"90",   x"29", 
  x"01",   x"B8",   x"B0",   x"09",   x"A0",   x"19",   x"11",   x"A8", 
  x"82",   x"3B",   x"33",   x"8A",   x"23",   x"9A",   x"92",   x"2B", 
  x"03",   x"BA",   x"B2",   x"0B",   x"A2",   x"1B",   x"13",   x"AA", 
  x"43",   x"FA",   x"F2",   x"4B",   x"E2",   x"5B",   x"53",   x"EA", 
  x"C2",   x"7B",   x"73",   x"CA",   x"63",   x"DA",   x"D2",   x"6B", 
  x"C3",   x"7A",   x"72",   x"CB",   x"62",   x"DB",   x"D3",   x"6A", 
  x"42",   x"FB",   x"F3",   x"4A",   x"E3",   x"5A",   x"52",   x"EB", 
  x"02",   x"BB",   x"B3",   x"0A",   x"A3",   x"1A",   x"12",   x"AB", 
  x"83",   x"3A",   x"32",   x"8B",   x"22",   x"9B",   x"93",   x"2A", 
  x"C7",   x"7E",   x"76",   x"CF",   x"66",   x"DF",   x"D7",   x"6E", 
  x"46",   x"FF",   x"F7",   x"4E",   x"E7",   x"5E",   x"56",   x"EF", 
  x"06",   x"BF",   x"B7",   x"0E",   x"A7",   x"1E",   x"16",   x"AF", 
  x"87",   x"3E",   x"36",   x"8F",   x"26",   x"9F",   x"97",   x"2E", 
  x"86",   x"3F",   x"37",   x"8E",   x"27",   x"9E",   x"96",   x"2F", 
  x"07",   x"BE",   x"B6",   x"0F",   x"A6",   x"1F",   x"17",   x"AE", 
  x"47",   x"FE",   x"F6",   x"4F",   x"E6",   x"5F",   x"57",   x"EE", 
  x"C6",   x"7F",   x"77",   x"CE",   x"67",   x"DE",   x"D6",   x"6F", 
  x"45",   x"FC",   x"F4",   x"4D",   x"E4",   x"5D",   x"55",   x"EC", 
  x"C4",   x"7D",   x"75",   x"CC",   x"65",   x"DC",   x"D4",   x"6D", 
  x"84",   x"3D",   x"35",   x"8C",   x"25",   x"9C",   x"94",   x"2D", 
  x"05",   x"BC",   x"B4",   x"0D",   x"A4",   x"1D",   x"15",   x"AC", 
  x"04",   x"BD",   x"B5",   x"0C",   x"A5",   x"1C",   x"14",   x"AD", 
  x"85",   x"3C",   x"34",   x"8D",   x"24",   x"9D",   x"95",   x"2C", 
  x"C5",   x"7C",   x"74",   x"CD",   x"64",   x"DD",   x"D5",   x"6C", 
  x"44",   x"FD",   x"F5",   x"4C",   x"E5",   x"5C",   x"54",   x"ED", 
  x"00",   x"BA",   x"B7",   x"0D",   x"AD",   x"17",   x"1A",   x"A0", 
  x"99",   x"23",   x"2E",   x"94",   x"34",   x"8E",   x"83",   x"39", 
  x"F1",   x"4B",   x"46",   x"FC",   x"5C",   x"E6",   x"EB",   x"51", 
  x"68",   x"D2",   x"DF",   x"65",   x"C5",   x"7F",   x"72",   x"C8", 
  x"21",   x"9B",   x"96",   x"2C",   x"8C",   x"36",   x"3B",   x"81", 
  x"B8",   x"02",   x"0F",   x"B5",   x"15",   x"AF",   x"A2",   x"18", 
  x"D0",   x"6A",   x"67",   x"DD",   x"7D",   x"C7",   x"CA",   x"70", 
  x"49",   x"F3",   x"FE",   x"44",   x"E4",   x"5E",   x"53",   x"E9", 
  x"42",   x"F8",   x"F5",   x"4F",   x"EF",   x"55",   x"58",   x"E2", 
  x"DB",   x"61",   x"6C",   x"D6",   x"76",   x"CC",   x"C1",   x"7B", 
  x"B3",   x"09",   x"04",   x"BE",   x"1E",   x"A4",   x"A9",   x"13", 
  x"2A",   x"90",   x"9D",   x"27",   x"87",   x"3D",   x"30",   x"8A", 
  x"63",   x"D9",   x"D4",   x"6E",   x"CE",   x"74",   x"79",   x"C3", 
  x"FA",   x"40",   x"4D",   x"F7",   x"57",   x"ED",   x"E0",   x"5A", 
  x"92",   x"28",   x"25",   x"9F",   x"3F",   x"85",   x"88",   x"32", 
  x"0B",   x"B1",   x"BC",   x"06",   x"A6",   x"1C",   x"11",   x"AB", 
  x"84",   x"3E",   x"33",   x"89",   x"29",   x"93",   x"9E",   x"24", 
  x"1D",   x"A7",   x"AA",   x"10",   x"B0",   x"0A",   x"07",   x"BD", 
  x"75",   x"CF",   x"C2",   x"78",   x"D8",   x"62",   x"6F",   x"D5", 
  x"EC",   x"56",   x"5B",   x"E1",   x"41",   x"FB",   x"F6",   x"4C", 
  x"A5",   x"1F",   x"12",   x"A8",   x"08",   x"B2",   x"BF",   x"05", 
  x"3C",   x"86",   x"8B",   x"31",   x"91",   x"2B",   x"26",   x"9C", 
  x"54",   x"EE",   x"E3",   x"59",   x"F9",   x"43",   x"4E",   x"F4", 
  x"CD",   x"77",   x"7A",   x"C0",   x"60",   x"DA",   x"D7",   x"6D", 
  x"C6",   x"7C",   x"71",   x"CB",   x"6B",   x"D1",   x"DC",   x"66", 
  x"5F",   x"E5",   x"E8",   x"52",   x"F2",   x"48",   x"45",   x"FF", 
  x"37",   x"8D",   x"80",   x"3A",   x"9A",   x"20",   x"2D",   x"97", 
  x"AE",   x"14",   x"19",   x"A3",   x"03",   x"B9",   x"B4",   x"0E", 
  x"E7",   x"5D",   x"50",   x"EA",   x"4A",   x"F0",   x"FD",   x"47", 
  x"7E",   x"C4",   x"C9",   x"73",   x"D3",   x"69",   x"64",   x"DE", 
  x"16",   x"AC",   x"A1",   x"1B",   x"BB",   x"01",   x"0C",   x"B6", 
  x"8F",   x"35",   x"38",   x"82",   x"22",   x"98",   x"95",   x"2F", 
  x"00",   x"BB",   x"B5",   x"0E",   x"A9",   x"12",   x"1C",   x"A7", 
  x"91",   x"2A",   x"24",   x"9F",   x"38",   x"83",   x"8D",   x"36", 
  x"E1",   x"5A",   x"54",   x"EF",   x"48",   x"F3",   x"FD",   x"46", 
  x"70",   x"CB",   x"C5",   x"7E",   x"D9",   x"62",   x"6C",   x"D7", 
  x"01",   x"BA",   x"B4",   x"0F",   x"A8",   x"13",   x"1D",   x"A6", 
  x"90",   x"2B",   x"25",   x"9E",   x"39",   x"82",   x"8C",   x"37", 
  x"E0",   x"5B",   x"55",   x"EE",   x"49",   x"F2",   x"FC",   x"47", 
  x"71",   x"CA",   x"C4",   x"7F",   x"D8",   x"63",   x"6D",   x"D6", 
  x"02",   x"B9",   x"B7",   x"0C",   x"AB",   x"10",   x"1E",   x"A5", 
  x"93",   x"28",   x"26",   x"9D",   x"3A",   x"81",   x"8F",   x"34", 
  x"E3",   x"58",   x"56",   x"ED",   x"4A",   x"F1",   x"FF",   x"44", 
  x"72",   x"C9",   x"C7",   x"7C",   x"DB",   x"60",   x"6E",   x"D5", 
  x"03",   x"B8",   x"B6",   x"0D",   x"AA",   x"11",   x"1F",   x"A4", 
  x"92",   x"29",   x"27",   x"9C",   x"3B",   x"80",   x"8E",   x"35", 
  x"E2",   x"59",   x"57",   x"EC",   x"4B",   x"F0",   x"FE",   x"45", 
  x"73",   x"C8",   x"C6",   x"7D",   x"DA",   x"61",   x"6F",   x"D4", 
  x"04",   x"BF",   x"B1",   x"0A",   x"AD",   x"16",   x"18",   x"A3", 
  x"95",   x"2E",   x"20",   x"9B",   x"3C",   x"87",   x"89",   x"32", 
  x"E5",   x"5E",   x"50",   x"EB",   x"4C",   x"F7",   x"F9",   x"42", 
  x"74",   x"CF",   x"C1",   x"7A",   x"DD",   x"66",   x"68",   x"D3", 
  x"05",   x"BE",   x"B0",   x"0B",   x"AC",   x"17",   x"19",   x"A2", 
  x"94",   x"2F",   x"21",   x"9A",   x"3D",   x"86",   x"88",   x"33", 
  x"E4",   x"5F",   x"51",   x"EA",   x"4D",   x"F6",   x"F8",   x"43", 
  x"75",   x"CE",   x"C0",   x"7B",   x"DC",   x"67",   x"69",   x"D2", 
  x"06",   x"BD",   x"B3",   x"08",   x"AF",   x"14",   x"1A",   x"A1", 
  x"97",   x"2C",   x"22",   x"99",   x"3E",   x"85",   x"8B",   x"30", 
  x"E7",   x"5C",   x"52",   x"E9",   x"4E",   x"F5",   x"FB",   x"40", 
  x"76",   x"CD",   x"C3",   x"78",   x"DF",   x"64",   x"6A",   x"D1", 
  x"07",   x"BC",   x"B2",   x"09",   x"AE",   x"15",   x"1B",   x"A0", 
  x"96",   x"2D",   x"23",   x"98",   x"3F",   x"84",   x"8A",   x"31", 
  x"E6",   x"5D",   x"53",   x"E8",   x"4F",   x"F4",   x"FA",   x"41", 
  x"77",   x"CC",   x"C2",   x"79",   x"DE",   x"65",   x"6B",   x"D0", 
  x"00",   x"BC",   x"BB",   x"07",   x"B5",   x"09",   x"0E",   x"B2", 
  x"A9",   x"15",   x"12",   x"AE",   x"1C",   x"A0",   x"A7",   x"1B", 
  x"91",   x"2D",   x"2A",   x"96",   x"24",   x"98",   x"9F",   x"23", 
  x"38",   x"84",   x"83",   x"3F",   x"8D",   x"31",   x"36",   x"8A", 
  x"E1",   x"5D",   x"5A",   x"E6",   x"54",   x"E8",   x"EF",   x"53", 
  x"48",   x"F4",   x"F3",   x"4F",   x"FD",   x"41",   x"46",   x"FA", 
  x"70",   x"CC",   x"CB",   x"77",   x"C5",   x"79",   x"7E",   x"C2", 
  x"D9",   x"65",   x"62",   x"DE",   x"6C",   x"D0",   x"D7",   x"6B", 
  x"01",   x"BD",   x"BA",   x"06",   x"B4",   x"08",   x"0F",   x"B3", 
  x"A8",   x"14",   x"13",   x"AF",   x"1D",   x"A1",   x"A6",   x"1A", 
  x"90",   x"2C",   x"2B",   x"97",   x"25",   x"99",   x"9E",   x"22", 
  x"39",   x"85",   x"82",   x"3E",   x"8C",   x"30",   x"37",   x"8B", 
  x"E0",   x"5C",   x"5B",   x"E7",   x"55",   x"E9",   x"EE",   x"52", 
  x"49",   x"F5",   x"F2",   x"4E",   x"FC",   x"40",   x"47",   x"FB", 
  x"71",   x"CD",   x"CA",   x"76",   x"C4",   x"78",   x"7F",   x"C3", 
  x"D8",   x"64",   x"63",   x"DF",   x"6D",   x"D1",   x"D6",   x"6A", 
  x"02",   x"BE",   x"B9",   x"05",   x"B7",   x"0B",   x"0C",   x"B0", 
  x"AB",   x"17",   x"10",   x"AC",   x"1E",   x"A2",   x"A5",   x"19", 
  x"93",   x"2F",   x"28",   x"94",   x"26",   x"9A",   x"9D",   x"21", 
  x"3A",   x"86",   x"81",   x"3D",   x"8F",   x"33",   x"34",   x"88", 
  x"E3",   x"5F",   x"58",   x"E4",   x"56",   x"EA",   x"ED",   x"51", 
  x"4A",   x"F6",   x"F1",   x"4D",   x"FF",   x"43",   x"44",   x"F8", 
  x"72",   x"CE",   x"C9",   x"75",   x"C7",   x"7B",   x"7C",   x"C0", 
  x"DB",   x"67",   x"60",   x"DC",   x"6E",   x"D2",   x"D5",   x"69", 
  x"03",   x"BF",   x"B8",   x"04",   x"B6",   x"0A",   x"0D",   x"B1", 
  x"AA",   x"16",   x"11",   x"AD",   x"1F",   x"A3",   x"A4",   x"18", 
  x"92",   x"2E",   x"29",   x"95",   x"27",   x"9B",   x"9C",   x"20", 
  x"3B",   x"87",   x"80",   x"3C",   x"8E",   x"32",   x"35",   x"89", 
  x"E2",   x"5E",   x"59",   x"E5",   x"57",   x"EB",   x"EC",   x"50", 
  x"4B",   x"F7",   x"F0",   x"4C",   x"FE",   x"42",   x"45",   x"F9", 
  x"73",   x"CF",   x"C8",   x"74",   x"C6",   x"7A",   x"7D",   x"C1", 
  x"DA",   x"66",   x"61",   x"DD",   x"6F",   x"D3",   x"D4",   x"68", 
  x"00",   x"BD",   x"B9",   x"04",   x"B1",   x"0C",   x"08",   x"B5", 
  x"A1",   x"1C",   x"18",   x"A5",   x"10",   x"AD",   x"A9",   x"14", 
  x"81",   x"3C",   x"38",   x"85",   x"30",   x"8D",   x"89",   x"34", 
  x"20",   x"9D",   x"99",   x"24",   x"91",   x"2C",   x"28",   x"95", 
  x"C1",   x"7C",   x"78",   x"C5",   x"70",   x"CD",   x"C9",   x"74", 
  x"60",   x"DD",   x"D9",   x"64",   x"D1",   x"6C",   x"68",   x"D5", 
  x"40",   x"FD",   x"F9",   x"44",   x"F1",   x"4C",   x"48",   x"F5", 
  x"E1",   x"5C",   x"58",   x"E5",   x"50",   x"ED",   x"E9",   x"54", 
  x"41",   x"FC",   x"F8",   x"45",   x"F0",   x"4D",   x"49",   x"F4", 
  x"E0",   x"5D",   x"59",   x"E4",   x"51",   x"EC",   x"E8",   x"55", 
  x"C0",   x"7D",   x"79",   x"C4",   x"71",   x"CC",   x"C8",   x"75", 
  x"61",   x"DC",   x"D8",   x"65",   x"D0",   x"6D",   x"69",   x"D4", 
  x"80",   x"3D",   x"39",   x"84",   x"31",   x"8C",   x"88",   x"35", 
  x"21",   x"9C",   x"98",   x"25",   x"90",   x"2D",   x"29",   x"94", 
  x"01",   x"BC",   x"B8",   x"05",   x"B0",   x"0D",   x"09",   x"B4", 
  x"A0",   x"1D",   x"19",   x"A4",   x"11",   x"AC",   x"A8",   x"15", 
  x"82",   x"3F",   x"3B",   x"86",   x"33",   x"8E",   x"8A",   x"37", 
  x"23",   x"9E",   x"9A",   x"27",   x"92",   x"2F",   x"2B",   x"96", 
  x"03",   x"BE",   x"BA",   x"07",   x"B2",   x"0F",   x"0B",   x"B6", 
  x"A2",   x"1F",   x"1B",   x"A6",   x"13",   x"AE",   x"AA",   x"17", 
  x"43",   x"FE",   x"FA",   x"47",   x"F2",   x"4F",   x"4B",   x"F6", 
  x"E2",   x"5F",   x"5B",   x"E6",   x"53",   x"EE",   x"EA",   x"57", 
  x"C2",   x"7F",   x"7B",   x"C6",   x"73",   x"CE",   x"CA",   x"77", 
  x"63",   x"DE",   x"DA",   x"67",   x"D2",   x"6F",   x"6B",   x"D6", 
  x"C3",   x"7E",   x"7A",   x"C7",   x"72",   x"CF",   x"CB",   x"76", 
  x"62",   x"DF",   x"DB",   x"66",   x"D3",   x"6E",   x"6A",   x"D7", 
  x"42",   x"FF",   x"FB",   x"46",   x"F3",   x"4E",   x"4A",   x"F7", 
  x"E3",   x"5E",   x"5A",   x"E7",   x"52",   x"EF",   x"EB",   x"56", 
  x"02",   x"BF",   x"BB",   x"06",   x"B3",   x"0E",   x"0A",   x"B7", 
  x"A3",   x"1E",   x"1A",   x"A7",   x"12",   x"AF",   x"AB",   x"16", 
  x"83",   x"3E",   x"3A",   x"87",   x"32",   x"8F",   x"8B",   x"36", 
  x"22",   x"9F",   x"9B",   x"26",   x"93",   x"2E",   x"2A",   x"97", 
  x"00",   x"BE",   x"BF",   x"01",   x"BD",   x"03",   x"02",   x"BC", 
  x"B9",   x"07",   x"06",   x"B8",   x"04",   x"BA",   x"BB",   x"05", 
  x"B1",   x"0F",   x"0E",   x"B0",   x"0C",   x"B2",   x"B3",   x"0D", 
  x"08",   x"B6",   x"B7",   x"09",   x"B5",   x"0B",   x"0A",   x"B4", 
  x"A1",   x"1F",   x"1E",   x"A0",   x"1C",   x"A2",   x"A3",   x"1D", 
  x"18",   x"A6",   x"A7",   x"19",   x"A5",   x"1B",   x"1A",   x"A4", 
  x"10",   x"AE",   x"AF",   x"11",   x"AD",   x"13",   x"12",   x"AC", 
  x"A9",   x"17",   x"16",   x"A8",   x"14",   x"AA",   x"AB",   x"15", 
  x"81",   x"3F",   x"3E",   x"80",   x"3C",   x"82",   x"83",   x"3D", 
  x"38",   x"86",   x"87",   x"39",   x"85",   x"3B",   x"3A",   x"84", 
  x"30",   x"8E",   x"8F",   x"31",   x"8D",   x"33",   x"32",   x"8C", 
  x"89",   x"37",   x"36",   x"88",   x"34",   x"8A",   x"8B",   x"35", 
  x"20",   x"9E",   x"9F",   x"21",   x"9D",   x"23",   x"22",   x"9C", 
  x"99",   x"27",   x"26",   x"98",   x"24",   x"9A",   x"9B",   x"25", 
  x"91",   x"2F",   x"2E",   x"90",   x"2C",   x"92",   x"93",   x"2D", 
  x"28",   x"96",   x"97",   x"29",   x"95",   x"2B",   x"2A",   x"94", 
  x"C1",   x"7F",   x"7E",   x"C0",   x"7C",   x"C2",   x"C3",   x"7D", 
  x"78",   x"C6",   x"C7",   x"79",   x"C5",   x"7B",   x"7A",   x"C4", 
  x"70",   x"CE",   x"CF",   x"71",   x"CD",   x"73",   x"72",   x"CC", 
  x"C9",   x"77",   x"76",   x"C8",   x"74",   x"CA",   x"CB",   x"75", 
  x"60",   x"DE",   x"DF",   x"61",   x"DD",   x"63",   x"62",   x"DC", 
  x"D9",   x"67",   x"66",   x"D8",   x"64",   x"DA",   x"DB",   x"65", 
  x"D1",   x"6F",   x"6E",   x"D0",   x"6C",   x"D2",   x"D3",   x"6D", 
  x"68",   x"D6",   x"D7",   x"69",   x"D5",   x"6B",   x"6A",   x"D4", 
  x"40",   x"FE",   x"FF",   x"41",   x"FD",   x"43",   x"42",   x"FC", 
  x"F9",   x"47",   x"46",   x"F8",   x"44",   x"FA",   x"FB",   x"45", 
  x"F1",   x"4F",   x"4E",   x"F0",   x"4C",   x"F2",   x"F3",   x"4D", 
  x"48",   x"F6",   x"F7",   x"49",   x"F5",   x"4B",   x"4A",   x"F4", 
  x"E1",   x"5F",   x"5E",   x"E0",   x"5C",   x"E2",   x"E3",   x"5D", 
  x"58",   x"E6",   x"E7",   x"59",   x"E5",   x"5B",   x"5A",   x"E4", 
  x"50",   x"EE",   x"EF",   x"51",   x"ED",   x"53",   x"52",   x"EC", 
  x"E9",   x"57",   x"56",   x"E8",   x"54",   x"EA",   x"EB",   x"55", 
  x"00",   x"BF",   x"BD",   x"02",   x"B9",   x"06",   x"04",   x"BB", 
  x"B1",   x"0E",   x"0C",   x"B3",   x"08",   x"B7",   x"B5",   x"0A", 
  x"A1",   x"1E",   x"1C",   x"A3",   x"18",   x"A7",   x"A5",   x"1A", 
  x"10",   x"AF",   x"AD",   x"12",   x"A9",   x"16",   x"14",   x"AB", 
  x"81",   x"3E",   x"3C",   x"83",   x"38",   x"87",   x"85",   x"3A", 
  x"30",   x"8F",   x"8D",   x"32",   x"89",   x"36",   x"34",   x"8B", 
  x"20",   x"9F",   x"9D",   x"22",   x"99",   x"26",   x"24",   x"9B", 
  x"91",   x"2E",   x"2C",   x"93",   x"28",   x"97",   x"95",   x"2A", 
  x"C1",   x"7E",   x"7C",   x"C3",   x"78",   x"C7",   x"C5",   x"7A", 
  x"70",   x"CF",   x"CD",   x"72",   x"C9",   x"76",   x"74",   x"CB", 
  x"60",   x"DF",   x"DD",   x"62",   x"D9",   x"66",   x"64",   x"DB", 
  x"D1",   x"6E",   x"6C",   x"D3",   x"68",   x"D7",   x"D5",   x"6A", 
  x"40",   x"FF",   x"FD",   x"42",   x"F9",   x"46",   x"44",   x"FB", 
  x"F1",   x"4E",   x"4C",   x"F3",   x"48",   x"F7",   x"F5",   x"4A", 
  x"E1",   x"5E",   x"5C",   x"E3",   x"58",   x"E7",   x"E5",   x"5A", 
  x"50",   x"EF",   x"ED",   x"52",   x"E9",   x"56",   x"54",   x"EB", 
  x"41",   x"FE",   x"FC",   x"43",   x"F8",   x"47",   x"45",   x"FA", 
  x"F0",   x"4F",   x"4D",   x"F2",   x"49",   x"F6",   x"F4",   x"4B", 
  x"E0",   x"5F",   x"5D",   x"E2",   x"59",   x"E6",   x"E4",   x"5B", 
  x"51",   x"EE",   x"EC",   x"53",   x"E8",   x"57",   x"55",   x"EA", 
  x"C0",   x"7F",   x"7D",   x"C2",   x"79",   x"C6",   x"C4",   x"7B", 
  x"71",   x"CE",   x"CC",   x"73",   x"C8",   x"77",   x"75",   x"CA", 
  x"61",   x"DE",   x"DC",   x"63",   x"D8",   x"67",   x"65",   x"DA", 
  x"D0",   x"6F",   x"6D",   x"D2",   x"69",   x"D6",   x"D4",   x"6B", 
  x"80",   x"3F",   x"3D",   x"82",   x"39",   x"86",   x"84",   x"3B", 
  x"31",   x"8E",   x"8C",   x"33",   x"88",   x"37",   x"35",   x"8A", 
  x"21",   x"9E",   x"9C",   x"23",   x"98",   x"27",   x"25",   x"9A", 
  x"90",   x"2F",   x"2D",   x"92",   x"29",   x"96",   x"94",   x"2B", 
  x"01",   x"BE",   x"BC",   x"03",   x"B8",   x"07",   x"05",   x"BA", 
  x"B0",   x"0F",   x"0D",   x"B2",   x"09",   x"B6",   x"B4",   x"0B", 
  x"A0",   x"1F",   x"1D",   x"A2",   x"19",   x"A6",   x"A4",   x"1B", 
  x"11",   x"AE",   x"AC",   x"13",   x"A8",   x"17",   x"15",   x"AA", 
  x"00",   x"C0",   x"43",   x"83",   x"86",   x"46",   x"C5",   x"05", 
  x"CF",   x"0F",   x"8C",   x"4C",   x"49",   x"89",   x"0A",   x"CA", 
  x"5D",   x"9D",   x"1E",   x"DE",   x"DB",   x"1B",   x"98",   x"58", 
  x"92",   x"52",   x"D1",   x"11",   x"14",   x"D4",   x"57",   x"97", 
  x"BA",   x"7A",   x"F9",   x"39",   x"3C",   x"FC",   x"7F",   x"BF", 
  x"75",   x"B5",   x"36",   x"F6",   x"F3",   x"33",   x"B0",   x"70", 
  x"E7",   x"27",   x"A4",   x"64",   x"61",   x"A1",   x"22",   x"E2", 
  x"28",   x"E8",   x"6B",   x"AB",   x"AE",   x"6E",   x"ED",   x"2D", 
  x"B7",   x"77",   x"F4",   x"34",   x"31",   x"F1",   x"72",   x"B2", 
  x"78",   x"B8",   x"3B",   x"FB",   x"FE",   x"3E",   x"BD",   x"7D", 
  x"EA",   x"2A",   x"A9",   x"69",   x"6C",   x"AC",   x"2F",   x"EF", 
  x"25",   x"E5",   x"66",   x"A6",   x"A3",   x"63",   x"E0",   x"20", 
  x"0D",   x"CD",   x"4E",   x"8E",   x"8B",   x"4B",   x"C8",   x"08", 
  x"C2",   x"02",   x"81",   x"41",   x"44",   x"84",   x"07",   x"C7", 
  x"50",   x"90",   x"13",   x"D3",   x"D6",   x"16",   x"95",   x"55", 
  x"9F",   x"5F",   x"DC",   x"1C",   x"19",   x"D9",   x"5A",   x"9A", 
  x"AD",   x"6D",   x"EE",   x"2E",   x"2B",   x"EB",   x"68",   x"A8", 
  x"62",   x"A2",   x"21",   x"E1",   x"E4",   x"24",   x"A7",   x"67", 
  x"F0",   x"30",   x"B3",   x"73",   x"76",   x"B6",   x"35",   x"F5", 
  x"3F",   x"FF",   x"7C",   x"BC",   x"B9",   x"79",   x"FA",   x"3A", 
  x"17",   x"D7",   x"54",   x"94",   x"91",   x"51",   x"D2",   x"12", 
  x"D8",   x"18",   x"9B",   x"5B",   x"5E",   x"9E",   x"1D",   x"DD", 
  x"4A",   x"8A",   x"09",   x"C9",   x"CC",   x"0C",   x"8F",   x"4F", 
  x"85",   x"45",   x"C6",   x"06",   x"03",   x"C3",   x"40",   x"80", 
  x"1A",   x"DA",   x"59",   x"99",   x"9C",   x"5C",   x"DF",   x"1F", 
  x"D5",   x"15",   x"96",   x"56",   x"53",   x"93",   x"10",   x"D0", 
  x"47",   x"87",   x"04",   x"C4",   x"C1",   x"01",   x"82",   x"42", 
  x"88",   x"48",   x"CB",   x"0B",   x"0E",   x"CE",   x"4D",   x"8D", 
  x"A0",   x"60",   x"E3",   x"23",   x"26",   x"E6",   x"65",   x"A5", 
  x"6F",   x"AF",   x"2C",   x"EC",   x"E9",   x"29",   x"AA",   x"6A", 
  x"FD",   x"3D",   x"BE",   x"7E",   x"7B",   x"BB",   x"38",   x"F8", 
  x"32",   x"F2",   x"71",   x"B1",   x"B4",   x"74",   x"F7",   x"37", 
  x"00",   x"C1",   x"41",   x"80",   x"82",   x"43",   x"C3",   x"02", 
  x"C7",   x"06",   x"86",   x"47",   x"45",   x"84",   x"04",   x"C5", 
  x"4D",   x"8C",   x"0C",   x"CD",   x"CF",   x"0E",   x"8E",   x"4F", 
  x"8A",   x"4B",   x"CB",   x"0A",   x"08",   x"C9",   x"49",   x"88", 
  x"9A",   x"5B",   x"DB",   x"1A",   x"18",   x"D9",   x"59",   x"98", 
  x"5D",   x"9C",   x"1C",   x"DD",   x"DF",   x"1E",   x"9E",   x"5F", 
  x"D7",   x"16",   x"96",   x"57",   x"55",   x"94",   x"14",   x"D5", 
  x"10",   x"D1",   x"51",   x"90",   x"92",   x"53",   x"D3",   x"12", 
  x"F7",   x"36",   x"B6",   x"77",   x"75",   x"B4",   x"34",   x"F5", 
  x"30",   x"F1",   x"71",   x"B0",   x"B2",   x"73",   x"F3",   x"32", 
  x"BA",   x"7B",   x"FB",   x"3A",   x"38",   x"F9",   x"79",   x"B8", 
  x"7D",   x"BC",   x"3C",   x"FD",   x"FF",   x"3E",   x"BE",   x"7F", 
  x"6D",   x"AC",   x"2C",   x"ED",   x"EF",   x"2E",   x"AE",   x"6F", 
  x"AA",   x"6B",   x"EB",   x"2A",   x"28",   x"E9",   x"69",   x"A8", 
  x"20",   x"E1",   x"61",   x"A0",   x"A2",   x"63",   x"E3",   x"22", 
  x"E7",   x"26",   x"A6",   x"67",   x"65",   x"A4",   x"24",   x"E5", 
  x"2D",   x"EC",   x"6C",   x"AD",   x"AF",   x"6E",   x"EE",   x"2F", 
  x"EA",   x"2B",   x"AB",   x"6A",   x"68",   x"A9",   x"29",   x"E8", 
  x"60",   x"A1",   x"21",   x"E0",   x"E2",   x"23",   x"A3",   x"62", 
  x"A7",   x"66",   x"E6",   x"27",   x"25",   x"E4",   x"64",   x"A5", 
  x"B7",   x"76",   x"F6",   x"37",   x"35",   x"F4",   x"74",   x"B5", 
  x"70",   x"B1",   x"31",   x"F0",   x"F2",   x"33",   x"B3",   x"72", 
  x"FA",   x"3B",   x"BB",   x"7A",   x"78",   x"B9",   x"39",   x"F8", 
  x"3D",   x"FC",   x"7C",   x"BD",   x"BF",   x"7E",   x"FE",   x"3F", 
  x"DA",   x"1B",   x"9B",   x"5A",   x"58",   x"99",   x"19",   x"D8", 
  x"1D",   x"DC",   x"5C",   x"9D",   x"9F",   x"5E",   x"DE",   x"1F", 
  x"97",   x"56",   x"D6",   x"17",   x"15",   x"D4",   x"54",   x"95", 
  x"50",   x"91",   x"11",   x"D0",   x"D2",   x"13",   x"93",   x"52", 
  x"40",   x"81",   x"01",   x"C0",   x"C2",   x"03",   x"83",   x"42", 
  x"87",   x"46",   x"C6",   x"07",   x"05",   x"C4",   x"44",   x"85", 
  x"0D",   x"CC",   x"4C",   x"8D",   x"8F",   x"4E",   x"CE",   x"0F", 
  x"CA",   x"0B",   x"8B",   x"4A",   x"48",   x"89",   x"09",   x"C8", 
  x"00",   x"C2",   x"47",   x"85",   x"8E",   x"4C",   x"C9",   x"0B", 
  x"DF",   x"1D",   x"98",   x"5A",   x"51",   x"93",   x"16",   x"D4", 
  x"7D",   x"BF",   x"3A",   x"F8",   x"F3",   x"31",   x"B4",   x"76", 
  x"A2",   x"60",   x"E5",   x"27",   x"2C",   x"EE",   x"6B",   x"A9", 
  x"FA",   x"38",   x"BD",   x"7F",   x"74",   x"B6",   x"33",   x"F1", 
  x"25",   x"E7",   x"62",   x"A0",   x"AB",   x"69",   x"EC",   x"2E", 
  x"87",   x"45",   x"C0",   x"02",   x"09",   x"CB",   x"4E",   x"8C", 
  x"58",   x"9A",   x"1F",   x"DD",   x"D6",   x"14",   x"91",   x"53", 
  x"37",   x"F5",   x"70",   x"B2",   x"B9",   x"7B",   x"FE",   x"3C", 
  x"E8",   x"2A",   x"AF",   x"6D",   x"66",   x"A4",   x"21",   x"E3", 
  x"4A",   x"88",   x"0D",   x"CF",   x"C4",   x"06",   x"83",   x"41", 
  x"95",   x"57",   x"D2",   x"10",   x"1B",   x"D9",   x"5C",   x"9E", 
  x"CD",   x"0F",   x"8A",   x"48",   x"43",   x"81",   x"04",   x"C6", 
  x"12",   x"D0",   x"55",   x"97",   x"9C",   x"5E",   x"DB",   x"19", 
  x"B0",   x"72",   x"F7",   x"35",   x"3E",   x"FC",   x"79",   x"BB", 
  x"6F",   x"AD",   x"28",   x"EA",   x"E1",   x"23",   x"A6",   x"64", 
  x"6E",   x"AC",   x"29",   x"EB",   x"E0",   x"22",   x"A7",   x"65", 
  x"B1",   x"73",   x"F6",   x"34",   x"3F",   x"FD",   x"78",   x"BA", 
  x"13",   x"D1",   x"54",   x"96",   x"9D",   x"5F",   x"DA",   x"18", 
  x"CC",   x"0E",   x"8B",   x"49",   x"42",   x"80",   x"05",   x"C7", 
  x"94",   x"56",   x"D3",   x"11",   x"1A",   x"D8",   x"5D",   x"9F", 
  x"4B",   x"89",   x"0C",   x"CE",   x"C5",   x"07",   x"82",   x"40", 
  x"E9",   x"2B",   x"AE",   x"6C",   x"67",   x"A5",   x"20",   x"E2", 
  x"36",   x"F4",   x"71",   x"B3",   x"B8",   x"7A",   x"FF",   x"3D", 
  x"59",   x"9B",   x"1E",   x"DC",   x"D7",   x"15",   x"90",   x"52", 
  x"86",   x"44",   x"C1",   x"03",   x"08",   x"CA",   x"4F",   x"8D", 
  x"24",   x"E6",   x"63",   x"A1",   x"AA",   x"68",   x"ED",   x"2F", 
  x"FB",   x"39",   x"BC",   x"7E",   x"75",   x"B7",   x"32",   x"F0", 
  x"A3",   x"61",   x"E4",   x"26",   x"2D",   x"EF",   x"6A",   x"A8", 
  x"7C",   x"BE",   x"3B",   x"F9",   x"F2",   x"30",   x"B5",   x"77", 
  x"DE",   x"1C",   x"99",   x"5B",   x"50",   x"92",   x"17",   x"D5", 
  x"01",   x"C3",   x"46",   x"84",   x"8F",   x"4D",   x"C8",   x"0A", 
  x"00",   x"C3",   x"45",   x"86",   x"8A",   x"49",   x"CF",   x"0C", 
  x"D7",   x"14",   x"92",   x"51",   x"5D",   x"9E",   x"18",   x"DB", 
  x"6D",   x"AE",   x"28",   x"EB",   x"E7",   x"24",   x"A2",   x"61", 
  x"BA",   x"79",   x"FF",   x"3C",   x"30",   x"F3",   x"75",   x"B6", 
  x"DA",   x"19",   x"9F",   x"5C",   x"50",   x"93",   x"15",   x"D6", 
  x"0D",   x"CE",   x"48",   x"8B",   x"87",   x"44",   x"C2",   x"01", 
  x"B7",   x"74",   x"F2",   x"31",   x"3D",   x"FE",   x"78",   x"BB", 
  x"60",   x"A3",   x"25",   x"E6",   x"EA",   x"29",   x"AF",   x"6C", 
  x"77",   x"B4",   x"32",   x"F1",   x"FD",   x"3E",   x"B8",   x"7B", 
  x"A0",   x"63",   x"E5",   x"26",   x"2A",   x"E9",   x"6F",   x"AC", 
  x"1A",   x"D9",   x"5F",   x"9C",   x"90",   x"53",   x"D5",   x"16", 
  x"CD",   x"0E",   x"88",   x"4B",   x"47",   x"84",   x"02",   x"C1", 
  x"AD",   x"6E",   x"E8",   x"2B",   x"27",   x"E4",   x"62",   x"A1", 
  x"7A",   x"B9",   x"3F",   x"FC",   x"F0",   x"33",   x"B5",   x"76", 
  x"C0",   x"03",   x"85",   x"46",   x"4A",   x"89",   x"0F",   x"CC", 
  x"17",   x"D4",   x"52",   x"91",   x"9D",   x"5E",   x"D8",   x"1B", 
  x"EE",   x"2D",   x"AB",   x"68",   x"64",   x"A7",   x"21",   x"E2", 
  x"39",   x"FA",   x"7C",   x"BF",   x"B3",   x"70",   x"F6",   x"35", 
  x"83",   x"40",   x"C6",   x"05",   x"09",   x"CA",   x"4C",   x"8F", 
  x"54",   x"97",   x"11",   x"D2",   x"DE",   x"1D",   x"9B",   x"58", 
  x"34",   x"F7",   x"71",   x"B2",   x"BE",   x"7D",   x"FB",   x"38", 
  x"E3",   x"20",   x"A6",   x"65",   x"69",   x"AA",   x"2C",   x"EF", 
  x"59",   x"9A",   x"1C",   x"DF",   x"D3",   x"10",   x"96",   x"55", 
  x"8E",   x"4D",   x"CB",   x"08",   x"04",   x"C7",   x"41",   x"82", 
  x"99",   x"5A",   x"DC",   x"1F",   x"13",   x"D0",   x"56",   x"95", 
  x"4E",   x"8D",   x"0B",   x"C8",   x"C4",   x"07",   x"81",   x"42", 
  x"F4",   x"37",   x"B1",   x"72",   x"7E",   x"BD",   x"3B",   x"F8", 
  x"23",   x"E0",   x"66",   x"A5",   x"A9",   x"6A",   x"EC",   x"2F", 
  x"43",   x"80",   x"06",   x"C5",   x"C9",   x"0A",   x"8C",   x"4F", 
  x"94",   x"57",   x"D1",   x"12",   x"1E",   x"DD",   x"5B",   x"98", 
  x"2E",   x"ED",   x"6B",   x"A8",   x"A4",   x"67",   x"E1",   x"22", 
  x"F9",   x"3A",   x"BC",   x"7F",   x"73",   x"B0",   x"36",   x"F5", 
  x"00",   x"C4",   x"4B",   x"8F",   x"96",   x"52",   x"DD",   x"19", 
  x"EF",   x"2B",   x"A4",   x"60",   x"79",   x"BD",   x"32",   x"F6", 
  x"1D",   x"D9",   x"56",   x"92",   x"8B",   x"4F",   x"C0",   x"04", 
  x"F2",   x"36",   x"B9",   x"7D",   x"64",   x"A0",   x"2F",   x"EB", 
  x"3A",   x"FE",   x"71",   x"B5",   x"AC",   x"68",   x"E7",   x"23", 
  x"D5",   x"11",   x"9E",   x"5A",   x"43",   x"87",   x"08",   x"CC", 
  x"27",   x"E3",   x"6C",   x"A8",   x"B1",   x"75",   x"FA",   x"3E", 
  x"C8",   x"0C",   x"83",   x"47",   x"5E",   x"9A",   x"15",   x"D1", 
  x"74",   x"B0",   x"3F",   x"FB",   x"E2",   x"26",   x"A9",   x"6D", 
  x"9B",   x"5F",   x"D0",   x"14",   x"0D",   x"C9",   x"46",   x"82", 
  x"69",   x"AD",   x"22",   x"E6",   x"FF",   x"3B",   x"B4",   x"70", 
  x"86",   x"42",   x"CD",   x"09",   x"10",   x"D4",   x"5B",   x"9F", 
  x"4E",   x"8A",   x"05",   x"C1",   x"D8",   x"1C",   x"93",   x"57", 
  x"A1",   x"65",   x"EA",   x"2E",   x"37",   x"F3",   x"7C",   x"B8", 
  x"53",   x"97",   x"18",   x"DC",   x"C5",   x"01",   x"8E",   x"4A", 
  x"BC",   x"78",   x"F7",   x"33",   x"2A",   x"EE",   x"61",   x"A5", 
  x"E8",   x"2C",   x"A3",   x"67",   x"7E",   x"BA",   x"35",   x"F1", 
  x"07",   x"C3",   x"4C",   x"88",   x"91",   x"55",   x"DA",   x"1E", 
  x"F5",   x"31",   x"BE",   x"7A",   x"63",   x"A7",   x"28",   x"EC", 
  x"1A",   x"DE",   x"51",   x"95",   x"8C",   x"48",   x"C7",   x"03", 
  x"D2",   x"16",   x"99",   x"5D",   x"44",   x"80",   x"0F",   x"CB", 
  x"3D",   x"F9",   x"76",   x"B2",   x"AB",   x"6F",   x"E0",   x"24", 
  x"CF",   x"0B",   x"84",   x"40",   x"59",   x"9D",   x"12",   x"D6", 
  x"20",   x"E4",   x"6B",   x"AF",   x"B6",   x"72",   x"FD",   x"39", 
  x"9C",   x"58",   x"D7",   x"13",   x"0A",   x"CE",   x"41",   x"85", 
  x"73",   x"B7",   x"38",   x"FC",   x"E5",   x"21",   x"AE",   x"6A", 
  x"81",   x"45",   x"CA",   x"0E",   x"17",   x"D3",   x"5C",   x"98", 
  x"6E",   x"AA",   x"25",   x"E1",   x"F8",   x"3C",   x"B3",   x"77", 
  x"A6",   x"62",   x"ED",   x"29",   x"30",   x"F4",   x"7B",   x"BF", 
  x"49",   x"8D",   x"02",   x"C6",   x"DF",   x"1B",   x"94",   x"50", 
  x"BB",   x"7F",   x"F0",   x"34",   x"2D",   x"E9",   x"66",   x"A2", 
  x"54",   x"90",   x"1F",   x"DB",   x"C2",   x"06",   x"89",   x"4D", 
  x"00",   x"C5",   x"49",   x"8C",   x"92",   x"57",   x"DB",   x"1E", 
  x"E7",   x"22",   x"AE",   x"6B",   x"75",   x"B0",   x"3C",   x"F9", 
  x"0D",   x"C8",   x"44",   x"81",   x"9F",   x"5A",   x"D6",   x"13", 
  x"EA",   x"2F",   x"A3",   x"66",   x"78",   x"BD",   x"31",   x"F4", 
  x"1A",   x"DF",   x"53",   x"96",   x"88",   x"4D",   x"C1",   x"04", 
  x"FD",   x"38",   x"B4",   x"71",   x"6F",   x"AA",   x"26",   x"E3", 
  x"17",   x"D2",   x"5E",   x"9B",   x"85",   x"40",   x"CC",   x"09", 
  x"F0",   x"35",   x"B9",   x"7C",   x"62",   x"A7",   x"2B",   x"EE", 
  x"34",   x"F1",   x"7D",   x"B8",   x"A6",   x"63",   x"EF",   x"2A", 
  x"D3",   x"16",   x"9A",   x"5F",   x"41",   x"84",   x"08",   x"CD", 
  x"39",   x"FC",   x"70",   x"B5",   x"AB",   x"6E",   x"E2",   x"27", 
  x"DE",   x"1B",   x"97",   x"52",   x"4C",   x"89",   x"05",   x"C0", 
  x"2E",   x"EB",   x"67",   x"A2",   x"BC",   x"79",   x"F5",   x"30", 
  x"C9",   x"0C",   x"80",   x"45",   x"5B",   x"9E",   x"12",   x"D7", 
  x"23",   x"E6",   x"6A",   x"AF",   x"B1",   x"74",   x"F8",   x"3D", 
  x"C4",   x"01",   x"8D",   x"48",   x"56",   x"93",   x"1F",   x"DA", 
  x"68",   x"AD",   x"21",   x"E4",   x"FA",   x"3F",   x"B3",   x"76", 
  x"8F",   x"4A",   x"C6",   x"03",   x"1D",   x"D8",   x"54",   x"91", 
  x"65",   x"A0",   x"2C",   x"E9",   x"F7",   x"32",   x"BE",   x"7B", 
  x"82",   x"47",   x"CB",   x"0E",   x"10",   x"D5",   x"59",   x"9C", 
  x"72",   x"B7",   x"3B",   x"FE",   x"E0",   x"25",   x"A9",   x"6C", 
  x"95",   x"50",   x"DC",   x"19",   x"07",   x"C2",   x"4E",   x"8B", 
  x"7F",   x"BA",   x"36",   x"F3",   x"ED",   x"28",   x"A4",   x"61", 
  x"98",   x"5D",   x"D1",   x"14",   x"0A",   x"CF",   x"43",   x"86", 
  x"5C",   x"99",   x"15",   x"D0",   x"CE",   x"0B",   x"87",   x"42", 
  x"BB",   x"7E",   x"F2",   x"37",   x"29",   x"EC",   x"60",   x"A5", 
  x"51",   x"94",   x"18",   x"DD",   x"C3",   x"06",   x"8A",   x"4F", 
  x"B6",   x"73",   x"FF",   x"3A",   x"24",   x"E1",   x"6D",   x"A8", 
  x"46",   x"83",   x"0F",   x"CA",   x"D4",   x"11",   x"9D",   x"58", 
  x"A1",   x"64",   x"E8",   x"2D",   x"33",   x"F6",   x"7A",   x"BF", 
  x"4B",   x"8E",   x"02",   x"C7",   x"D9",   x"1C",   x"90",   x"55", 
  x"AC",   x"69",   x"E5",   x"20",   x"3E",   x"FB",   x"77",   x"B2", 
  x"00",   x"C6",   x"4F",   x"89",   x"9E",   x"58",   x"D1",   x"17", 
  x"FF",   x"39",   x"B0",   x"76",   x"61",   x"A7",   x"2E",   x"E8", 
  x"3D",   x"FB",   x"72",   x"B4",   x"A3",   x"65",   x"EC",   x"2A", 
  x"C2",   x"04",   x"8D",   x"4B",   x"5C",   x"9A",   x"13",   x"D5", 
  x"7A",   x"BC",   x"35",   x"F3",   x"E4",   x"22",   x"AB",   x"6D", 
  x"85",   x"43",   x"CA",   x"0C",   x"1B",   x"DD",   x"54",   x"92", 
  x"47",   x"81",   x"08",   x"CE",   x"D9",   x"1F",   x"96",   x"50", 
  x"B8",   x"7E",   x"F7",   x"31",   x"26",   x"E0",   x"69",   x"AF", 
  x"F4",   x"32",   x"BB",   x"7D",   x"6A",   x"AC",   x"25",   x"E3", 
  x"0B",   x"CD",   x"44",   x"82",   x"95",   x"53",   x"DA",   x"1C", 
  x"C9",   x"0F",   x"86",   x"40",   x"57",   x"91",   x"18",   x"DE", 
  x"36",   x"F0",   x"79",   x"BF",   x"A8",   x"6E",   x"E7",   x"21", 
  x"8E",   x"48",   x"C1",   x"07",   x"10",   x"D6",   x"5F",   x"99", 
  x"71",   x"B7",   x"3E",   x"F8",   x"EF",   x"29",   x"A0",   x"66", 
  x"B3",   x"75",   x"FC",   x"3A",   x"2D",   x"EB",   x"62",   x"A4", 
  x"4C",   x"8A",   x"03",   x"C5",   x"D2",   x"14",   x"9D",   x"5B", 
  x"2B",   x"ED",   x"64",   x"A2",   x"B5",   x"73",   x"FA",   x"3C", 
  x"D4",   x"12",   x"9B",   x"5D",   x"4A",   x"8C",   x"05",   x"C3", 
  x"16",   x"D0",   x"59",   x"9F",   x"88",   x"4E",   x"C7",   x"01", 
  x"E9",   x"2F",   x"A6",   x"60",   x"77",   x"B1",   x"38",   x"FE", 
  x"51",   x"97",   x"1E",   x"D8",   x"CF",   x"09",   x"80",   x"46", 
  x"AE",   x"68",   x"E1",   x"27",   x"30",   x"F6",   x"7F",   x"B9", 
  x"6C",   x"AA",   x"23",   x"E5",   x"F2",   x"34",   x"BD",   x"7B", 
  x"93",   x"55",   x"DC",   x"1A",   x"0D",   x"CB",   x"42",   x"84", 
  x"DF",   x"19",   x"90",   x"56",   x"41",   x"87",   x"0E",   x"C8", 
  x"20",   x"E6",   x"6F",   x"A9",   x"BE",   x"78",   x"F1",   x"37", 
  x"E2",   x"24",   x"AD",   x"6B",   x"7C",   x"BA",   x"33",   x"F5", 
  x"1D",   x"DB",   x"52",   x"94",   x"83",   x"45",   x"CC",   x"0A", 
  x"A5",   x"63",   x"EA",   x"2C",   x"3B",   x"FD",   x"74",   x"B2", 
  x"5A",   x"9C",   x"15",   x"D3",   x"C4",   x"02",   x"8B",   x"4D", 
  x"98",   x"5E",   x"D7",   x"11",   x"06",   x"C0",   x"49",   x"8F", 
  x"67",   x"A1",   x"28",   x"EE",   x"F9",   x"3F",   x"B6",   x"70", 
  x"00",   x"C7",   x"4D",   x"8A",   x"9A",   x"5D",   x"D7",   x"10", 
  x"F7",   x"30",   x"BA",   x"7D",   x"6D",   x"AA",   x"20",   x"E7", 
  x"2D",   x"EA",   x"60",   x"A7",   x"B7",   x"70",   x"FA",   x"3D", 
  x"DA",   x"1D",   x"97",   x"50",   x"40",   x"87",   x"0D",   x"CA", 
  x"5A",   x"9D",   x"17",   x"D0",   x"C0",   x"07",   x"8D",   x"4A", 
  x"AD",   x"6A",   x"E0",   x"27",   x"37",   x"F0",   x"7A",   x"BD", 
  x"77",   x"B0",   x"3A",   x"FD",   x"ED",   x"2A",   x"A0",   x"67", 
  x"80",   x"47",   x"CD",   x"0A",   x"1A",   x"DD",   x"57",   x"90", 
  x"B4",   x"73",   x"F9",   x"3E",   x"2E",   x"E9",   x"63",   x"A4", 
  x"43",   x"84",   x"0E",   x"C9",   x"D9",   x"1E",   x"94",   x"53", 
  x"99",   x"5E",   x"D4",   x"13",   x"03",   x"C4",   x"4E",   x"89", 
  x"6E",   x"A9",   x"23",   x"E4",   x"F4",   x"33",   x"B9",   x"7E", 
  x"EE",   x"29",   x"A3",   x"64",   x"74",   x"B3",   x"39",   x"FE", 
  x"19",   x"DE",   x"54",   x"93",   x"83",   x"44",   x"CE",   x"09", 
  x"C3",   x"04",   x"8E",   x"49",   x"59",   x"9E",   x"14",   x"D3", 
  x"34",   x"F3",   x"79",   x"BE",   x"AE",   x"69",   x"E3",   x"24", 
  x"AB",   x"6C",   x"E6",   x"21",   x"31",   x"F6",   x"7C",   x"BB", 
  x"5C",   x"9B",   x"11",   x"D6",   x"C6",   x"01",   x"8B",   x"4C", 
  x"86",   x"41",   x"CB",   x"0C",   x"1C",   x"DB",   x"51",   x"96", 
  x"71",   x"B6",   x"3C",   x"FB",   x"EB",   x"2C",   x"A6",   x"61", 
  x"F1",   x"36",   x"BC",   x"7B",   x"6B",   x"AC",   x"26",   x"E1", 
  x"06",   x"C1",   x"4B",   x"8C",   x"9C",   x"5B",   x"D1",   x"16", 
  x"DC",   x"1B",   x"91",   x"56",   x"46",   x"81",   x"0B",   x"CC", 
  x"2B",   x"EC",   x"66",   x"A1",   x"B1",   x"76",   x"FC",   x"3B", 
  x"1F",   x"D8",   x"52",   x"95",   x"85",   x"42",   x"C8",   x"0F", 
  x"E8",   x"2F",   x"A5",   x"62",   x"72",   x"B5",   x"3F",   x"F8", 
  x"32",   x"F5",   x"7F",   x"B8",   x"A8",   x"6F",   x"E5",   x"22", 
  x"C5",   x"02",   x"88",   x"4F",   x"5F",   x"98",   x"12",   x"D5", 
  x"45",   x"82",   x"08",   x"CF",   x"DF",   x"18",   x"92",   x"55", 
  x"B2",   x"75",   x"FF",   x"38",   x"28",   x"EF",   x"65",   x"A2", 
  x"68",   x"AF",   x"25",   x"E2",   x"F2",   x"35",   x"BF",   x"78", 
  x"9F",   x"58",   x"D2",   x"15",   x"05",   x"C2",   x"48",   x"8F", 
  x"00",   x"C8",   x"53",   x"9B",   x"A6",   x"6E",   x"F5",   x"3D", 
  x"8F",   x"47",   x"DC",   x"14",   x"29",   x"E1",   x"7A",   x"B2", 
  x"DD",   x"15",   x"8E",   x"46",   x"7B",   x"B3",   x"28",   x"E0", 
  x"52",   x"9A",   x"01",   x"C9",   x"F4",   x"3C",   x"A7",   x"6F", 
  x"79",   x"B1",   x"2A",   x"E2",   x"DF",   x"17",   x"8C",   x"44", 
  x"F6",   x"3E",   x"A5",   x"6D",   x"50",   x"98",   x"03",   x"CB", 
  x"A4",   x"6C",   x"F7",   x"3F",   x"02",   x"CA",   x"51",   x"99", 
  x"2B",   x"E3",   x"78",   x"B0",   x"8D",   x"45",   x"DE",   x"16", 
  x"F2",   x"3A",   x"A1",   x"69",   x"54",   x"9C",   x"07",   x"CF", 
  x"7D",   x"B5",   x"2E",   x"E6",   x"DB",   x"13",   x"88",   x"40", 
  x"2F",   x"E7",   x"7C",   x"B4",   x"89",   x"41",   x"DA",   x"12", 
  x"A0",   x"68",   x"F3",   x"3B",   x"06",   x"CE",   x"55",   x"9D", 
  x"8B",   x"43",   x"D8",   x"10",   x"2D",   x"E5",   x"7E",   x"B6", 
  x"04",   x"CC",   x"57",   x"9F",   x"A2",   x"6A",   x"F1",   x"39", 
  x"56",   x"9E",   x"05",   x"CD",   x"F0",   x"38",   x"A3",   x"6B", 
  x"D9",   x"11",   x"8A",   x"42",   x"7F",   x"B7",   x"2C",   x"E4", 
  x"27",   x"EF",   x"74",   x"BC",   x"81",   x"49",   x"D2",   x"1A", 
  x"A8",   x"60",   x"FB",   x"33",   x"0E",   x"C6",   x"5D",   x"95", 
  x"FA",   x"32",   x"A9",   x"61",   x"5C",   x"94",   x"0F",   x"C7", 
  x"75",   x"BD",   x"26",   x"EE",   x"D3",   x"1B",   x"80",   x"48", 
  x"5E",   x"96",   x"0D",   x"C5",   x"F8",   x"30",   x"AB",   x"63", 
  x"D1",   x"19",   x"82",   x"4A",   x"77",   x"BF",   x"24",   x"EC", 
  x"83",   x"4B",   x"D0",   x"18",   x"25",   x"ED",   x"76",   x"BE", 
  x"0C",   x"C4",   x"5F",   x"97",   x"AA",   x"62",   x"F9",   x"31", 
  x"D5",   x"1D",   x"86",   x"4E",   x"73",   x"BB",   x"20",   x"E8", 
  x"5A",   x"92",   x"09",   x"C1",   x"FC",   x"34",   x"AF",   x"67", 
  x"08",   x"C0",   x"5B",   x"93",   x"AE",   x"66",   x"FD",   x"35", 
  x"87",   x"4F",   x"D4",   x"1C",   x"21",   x"E9",   x"72",   x"BA", 
  x"AC",   x"64",   x"FF",   x"37",   x"0A",   x"C2",   x"59",   x"91", 
  x"23",   x"EB",   x"70",   x"B8",   x"85",   x"4D",   x"D6",   x"1E", 
  x"71",   x"B9",   x"22",   x"EA",   x"D7",   x"1F",   x"84",   x"4C", 
  x"FE",   x"36",   x"AD",   x"65",   x"58",   x"90",   x"0B",   x"C3", 
  x"00",   x"C9",   x"51",   x"98",   x"A2",   x"6B",   x"F3",   x"3A", 
  x"87",   x"4E",   x"D6",   x"1F",   x"25",   x"EC",   x"74",   x"BD", 
  x"CD",   x"04",   x"9C",   x"55",   x"6F",   x"A6",   x"3E",   x"F7", 
  x"4A",   x"83",   x"1B",   x"D2",   x"E8",   x"21",   x"B9",   x"70", 
  x"59",   x"90",   x"08",   x"C1",   x"FB",   x"32",   x"AA",   x"63", 
  x"DE",   x"17",   x"8F",   x"46",   x"7C",   x"B5",   x"2D",   x"E4", 
  x"94",   x"5D",   x"C5",   x"0C",   x"36",   x"FF",   x"67",   x"AE", 
  x"13",   x"DA",   x"42",   x"8B",   x"B1",   x"78",   x"E0",   x"29", 
  x"B2",   x"7B",   x"E3",   x"2A",   x"10",   x"D9",   x"41",   x"88", 
  x"35",   x"FC",   x"64",   x"AD",   x"97",   x"5E",   x"C6",   x"0F", 
  x"7F",   x"B6",   x"2E",   x"E7",   x"DD",   x"14",   x"8C",   x"45", 
  x"F8",   x"31",   x"A9",   x"60",   x"5A",   x"93",   x"0B",   x"C2", 
  x"EB",   x"22",   x"BA",   x"73",   x"49",   x"80",   x"18",   x"D1", 
  x"6C",   x"A5",   x"3D",   x"F4",   x"CE",   x"07",   x"9F",   x"56", 
  x"26",   x"EF",   x"77",   x"BE",   x"84",   x"4D",   x"D5",   x"1C", 
  x"A1",   x"68",   x"F0",   x"39",   x"03",   x"CA",   x"52",   x"9B", 
  x"A7",   x"6E",   x"F6",   x"3F",   x"05",   x"CC",   x"54",   x"9D", 
  x"20",   x"E9",   x"71",   x"B8",   x"82",   x"4B",   x"D3",   x"1A", 
  x"6A",   x"A3",   x"3B",   x"F2",   x"C8",   x"01",   x"99",   x"50", 
  x"ED",   x"24",   x"BC",   x"75",   x"4F",   x"86",   x"1E",   x"D7", 
  x"FE",   x"37",   x"AF",   x"66",   x"5C",   x"95",   x"0D",   x"C4", 
  x"79",   x"B0",   x"28",   x"E1",   x"DB",   x"12",   x"8A",   x"43", 
  x"33",   x"FA",   x"62",   x"AB",   x"91",   x"58",   x"C0",   x"09", 
  x"B4",   x"7D",   x"E5",   x"2C",   x"16",   x"DF",   x"47",   x"8E", 
  x"15",   x"DC",   x"44",   x"8D",   x"B7",   x"7E",   x"E6",   x"2F", 
  x"92",   x"5B",   x"C3",   x"0A",   x"30",   x"F9",   x"61",   x"A8", 
  x"D8",   x"11",   x"89",   x"40",   x"7A",   x"B3",   x"2B",   x"E2", 
  x"5F",   x"96",   x"0E",   x"C7",   x"FD",   x"34",   x"AC",   x"65", 
  x"4C",   x"85",   x"1D",   x"D4",   x"EE",   x"27",   x"BF",   x"76", 
  x"CB",   x"02",   x"9A",   x"53",   x"69",   x"A0",   x"38",   x"F1", 
  x"81",   x"48",   x"D0",   x"19",   x"23",   x"EA",   x"72",   x"BB", 
  x"06",   x"CF",   x"57",   x"9E",   x"A4",   x"6D",   x"F5",   x"3C", 
  x"00",   x"CA",   x"57",   x"9D",   x"AE",   x"64",   x"F9",   x"33", 
  x"9F",   x"55",   x"C8",   x"02",   x"31",   x"FB",   x"66",   x"AC", 
  x"FD",   x"37",   x"AA",   x"60",   x"53",   x"99",   x"04",   x"CE", 
  x"62",   x"A8",   x"35",   x"FF",   x"CC",   x"06",   x"9B",   x"51", 
  x"39",   x"F3",   x"6E",   x"A4",   x"97",   x"5D",   x"C0",   x"0A", 
  x"A6",   x"6C",   x"F1",   x"3B",   x"08",   x"C2",   x"5F",   x"95", 
  x"C4",   x"0E",   x"93",   x"59",   x"6A",   x"A0",   x"3D",   x"F7", 
  x"5B",   x"91",   x"0C",   x"C6",   x"F5",   x"3F",   x"A2",   x"68", 
  x"72",   x"B8",   x"25",   x"EF",   x"DC",   x"16",   x"8B",   x"41", 
  x"ED",   x"27",   x"BA",   x"70",   x"43",   x"89",   x"14",   x"DE", 
  x"8F",   x"45",   x"D8",   x"12",   x"21",   x"EB",   x"76",   x"BC", 
  x"10",   x"DA",   x"47",   x"8D",   x"BE",   x"74",   x"E9",   x"23", 
  x"4B",   x"81",   x"1C",   x"D6",   x"E5",   x"2F",   x"B2",   x"78", 
  x"D4",   x"1E",   x"83",   x"49",   x"7A",   x"B0",   x"2D",   x"E7", 
  x"B6",   x"7C",   x"E1",   x"2B",   x"18",   x"D2",   x"4F",   x"85", 
  x"29",   x"E3",   x"7E",   x"B4",   x"87",   x"4D",   x"D0",   x"1A", 
  x"E4",   x"2E",   x"B3",   x"79",   x"4A",   x"80",   x"1D",   x"D7", 
  x"7B",   x"B1",   x"2C",   x"E6",   x"D5",   x"1F",   x"82",   x"48", 
  x"19",   x"D3",   x"4E",   x"84",   x"B7",   x"7D",   x"E0",   x"2A", 
  x"86",   x"4C",   x"D1",   x"1B",   x"28",   x"E2",   x"7F",   x"B5", 
  x"DD",   x"17",   x"8A",   x"40",   x"73",   x"B9",   x"24",   x"EE", 
  x"42",   x"88",   x"15",   x"DF",   x"EC",   x"26",   x"BB",   x"71", 
  x"20",   x"EA",   x"77",   x"BD",   x"8E",   x"44",   x"D9",   x"13", 
  x"BF",   x"75",   x"E8",   x"22",   x"11",   x"DB",   x"46",   x"8C", 
  x"96",   x"5C",   x"C1",   x"0B",   x"38",   x"F2",   x"6F",   x"A5", 
  x"09",   x"C3",   x"5E",   x"94",   x"A7",   x"6D",   x"F0",   x"3A", 
  x"6B",   x"A1",   x"3C",   x"F6",   x"C5",   x"0F",   x"92",   x"58", 
  x"F4",   x"3E",   x"A3",   x"69",   x"5A",   x"90",   x"0D",   x"C7", 
  x"AF",   x"65",   x"F8",   x"32",   x"01",   x"CB",   x"56",   x"9C", 
  x"30",   x"FA",   x"67",   x"AD",   x"9E",   x"54",   x"C9",   x"03", 
  x"52",   x"98",   x"05",   x"CF",   x"FC",   x"36",   x"AB",   x"61", 
  x"CD",   x"07",   x"9A",   x"50",   x"63",   x"A9",   x"34",   x"FE", 
  x"00",   x"CB",   x"55",   x"9E",   x"AA",   x"61",   x"FF",   x"34", 
  x"97",   x"5C",   x"C2",   x"09",   x"3D",   x"F6",   x"68",   x"A3", 
  x"ED",   x"26",   x"B8",   x"73",   x"47",   x"8C",   x"12",   x"D9", 
  x"7A",   x"B1",   x"2F",   x"E4",   x"D0",   x"1B",   x"85",   x"4E", 
  x"19",   x"D2",   x"4C",   x"87",   x"B3",   x"78",   x"E6",   x"2D", 
  x"8E",   x"45",   x"DB",   x"10",   x"24",   x"EF",   x"71",   x"BA", 
  x"F4",   x"3F",   x"A1",   x"6A",   x"5E",   x"95",   x"0B",   x"C0", 
  x"63",   x"A8",   x"36",   x"FD",   x"C9",   x"02",   x"9C",   x"57", 
  x"32",   x"F9",   x"67",   x"AC",   x"98",   x"53",   x"CD",   x"06", 
  x"A5",   x"6E",   x"F0",   x"3B",   x"0F",   x"C4",   x"5A",   x"91", 
  x"DF",   x"14",   x"8A",   x"41",   x"75",   x"BE",   x"20",   x"EB", 
  x"48",   x"83",   x"1D",   x"D6",   x"E2",   x"29",   x"B7",   x"7C", 
  x"2B",   x"E0",   x"7E",   x"B5",   x"81",   x"4A",   x"D4",   x"1F", 
  x"BC",   x"77",   x"E9",   x"22",   x"16",   x"DD",   x"43",   x"88", 
  x"C6",   x"0D",   x"93",   x"58",   x"6C",   x"A7",   x"39",   x"F2", 
  x"51",   x"9A",   x"04",   x"CF",   x"FB",   x"30",   x"AE",   x"65", 
  x"64",   x"AF",   x"31",   x"FA",   x"CE",   x"05",   x"9B",   x"50", 
  x"F3",   x"38",   x"A6",   x"6D",   x"59",   x"92",   x"0C",   x"C7", 
  x"89",   x"42",   x"DC",   x"17",   x"23",   x"E8",   x"76",   x"BD", 
  x"1E",   x"D5",   x"4B",   x"80",   x"B4",   x"7F",   x"E1",   x"2A", 
  x"7D",   x"B6",   x"28",   x"E3",   x"D7",   x"1C",   x"82",   x"49", 
  x"EA",   x"21",   x"BF",   x"74",   x"40",   x"8B",   x"15",   x"DE", 
  x"90",   x"5B",   x"C5",   x"0E",   x"3A",   x"F1",   x"6F",   x"A4", 
  x"07",   x"CC",   x"52",   x"99",   x"AD",   x"66",   x"F8",   x"33", 
  x"56",   x"9D",   x"03",   x"C8",   x"FC",   x"37",   x"A9",   x"62", 
  x"C1",   x"0A",   x"94",   x"5F",   x"6B",   x"A0",   x"3E",   x"F5", 
  x"BB",   x"70",   x"EE",   x"25",   x"11",   x"DA",   x"44",   x"8F", 
  x"2C",   x"E7",   x"79",   x"B2",   x"86",   x"4D",   x"D3",   x"18", 
  x"4F",   x"84",   x"1A",   x"D1",   x"E5",   x"2E",   x"B0",   x"7B", 
  x"D8",   x"13",   x"8D",   x"46",   x"72",   x"B9",   x"27",   x"EC", 
  x"A2",   x"69",   x"F7",   x"3C",   x"08",   x"C3",   x"5D",   x"96", 
  x"35",   x"FE",   x"60",   x"AB",   x"9F",   x"54",   x"CA",   x"01", 
  x"00",   x"CC",   x"5B",   x"97",   x"B6",   x"7A",   x"ED",   x"21", 
  x"AF",   x"63",   x"F4",   x"38",   x"19",   x"D5",   x"42",   x"8E", 
  x"9D",   x"51",   x"C6",   x"0A",   x"2B",   x"E7",   x"70",   x"BC", 
  x"32",   x"FE",   x"69",   x"A5",   x"84",   x"48",   x"DF",   x"13", 
  x"F9",   x"35",   x"A2",   x"6E",   x"4F",   x"83",   x"14",   x"D8", 
  x"56",   x"9A",   x"0D",   x"C1",   x"E0",   x"2C",   x"BB",   x"77", 
  x"64",   x"A8",   x"3F",   x"F3",   x"D2",   x"1E",   x"89",   x"45", 
  x"CB",   x"07",   x"90",   x"5C",   x"7D",   x"B1",   x"26",   x"EA", 
  x"31",   x"FD",   x"6A",   x"A6",   x"87",   x"4B",   x"DC",   x"10", 
  x"9E",   x"52",   x"C5",   x"09",   x"28",   x"E4",   x"73",   x"BF", 
  x"AC",   x"60",   x"F7",   x"3B",   x"1A",   x"D6",   x"41",   x"8D", 
  x"03",   x"CF",   x"58",   x"94",   x"B5",   x"79",   x"EE",   x"22", 
  x"C8",   x"04",   x"93",   x"5F",   x"7E",   x"B2",   x"25",   x"E9", 
  x"67",   x"AB",   x"3C",   x"F0",   x"D1",   x"1D",   x"8A",   x"46", 
  x"55",   x"99",   x"0E",   x"C2",   x"E3",   x"2F",   x"B8",   x"74", 
  x"FA",   x"36",   x"A1",   x"6D",   x"4C",   x"80",   x"17",   x"DB", 
  x"62",   x"AE",   x"39",   x"F5",   x"D4",   x"18",   x"8F",   x"43", 
  x"CD",   x"01",   x"96",   x"5A",   x"7B",   x"B7",   x"20",   x"EC", 
  x"FF",   x"33",   x"A4",   x"68",   x"49",   x"85",   x"12",   x"DE", 
  x"50",   x"9C",   x"0B",   x"C7",   x"E6",   x"2A",   x"BD",   x"71", 
  x"9B",   x"57",   x"C0",   x"0C",   x"2D",   x"E1",   x"76",   x"BA", 
  x"34",   x"F8",   x"6F",   x"A3",   x"82",   x"4E",   x"D9",   x"15", 
  x"06",   x"CA",   x"5D",   x"91",   x"B0",   x"7C",   x"EB",   x"27", 
  x"A9",   x"65",   x"F2",   x"3E",   x"1F",   x"D3",   x"44",   x"88", 
  x"53",   x"9F",   x"08",   x"C4",   x"E5",   x"29",   x"BE",   x"72", 
  x"FC",   x"30",   x"A7",   x"6B",   x"4A",   x"86",   x"11",   x"DD", 
  x"CE",   x"02",   x"95",   x"59",   x"78",   x"B4",   x"23",   x"EF", 
  x"61",   x"AD",   x"3A",   x"F6",   x"D7",   x"1B",   x"8C",   x"40", 
  x"AA",   x"66",   x"F1",   x"3D",   x"1C",   x"D0",   x"47",   x"8B", 
  x"05",   x"C9",   x"5E",   x"92",   x"B3",   x"7F",   x"E8",   x"24", 
  x"37",   x"FB",   x"6C",   x"A0",   x"81",   x"4D",   x"DA",   x"16", 
  x"98",   x"54",   x"C3",   x"0F",   x"2E",   x"E2",   x"75",   x"B9", 
  x"00",   x"CD",   x"59",   x"94",   x"B2",   x"7F",   x"EB",   x"26", 
  x"A7",   x"6A",   x"FE",   x"33",   x"15",   x"D8",   x"4C",   x"81", 
  x"8D",   x"40",   x"D4",   x"19",   x"3F",   x"F2",   x"66",   x"AB", 
  x"2A",   x"E7",   x"73",   x"BE",   x"98",   x"55",   x"C1",   x"0C", 
  x"D9",   x"14",   x"80",   x"4D",   x"6B",   x"A6",   x"32",   x"FF", 
  x"7E",   x"B3",   x"27",   x"EA",   x"CC",   x"01",   x"95",   x"58", 
  x"54",   x"99",   x"0D",   x"C0",   x"E6",   x"2B",   x"BF",   x"72", 
  x"F3",   x"3E",   x"AA",   x"67",   x"41",   x"8C",   x"18",   x"D5", 
  x"71",   x"BC",   x"28",   x"E5",   x"C3",   x"0E",   x"9A",   x"57", 
  x"D6",   x"1B",   x"8F",   x"42",   x"64",   x"A9",   x"3D",   x"F0", 
  x"FC",   x"31",   x"A5",   x"68",   x"4E",   x"83",   x"17",   x"DA", 
  x"5B",   x"96",   x"02",   x"CF",   x"E9",   x"24",   x"B0",   x"7D", 
  x"A8",   x"65",   x"F1",   x"3C",   x"1A",   x"D7",   x"43",   x"8E", 
  x"0F",   x"C2",   x"56",   x"9B",   x"BD",   x"70",   x"E4",   x"29", 
  x"25",   x"E8",   x"7C",   x"B1",   x"97",   x"5A",   x"CE",   x"03", 
  x"82",   x"4F",   x"DB",   x"16",   x"30",   x"FD",   x"69",   x"A4", 
  x"E2",   x"2F",   x"BB",   x"76",   x"50",   x"9D",   x"09",   x"C4", 
  x"45",   x"88",   x"1C",   x"D1",   x"F7",   x"3A",   x"AE",   x"63", 
  x"6F",   x"A2",   x"36",   x"FB",   x"DD",   x"10",   x"84",   x"49", 
  x"C8",   x"05",   x"91",   x"5C",   x"7A",   x"B7",   x"23",   x"EE", 
  x"3B",   x"F6",   x"62",   x"AF",   x"89",   x"44",   x"D0",   x"1D", 
  x"9C",   x"51",   x"C5",   x"08",   x"2E",   x"E3",   x"77",   x"BA", 
  x"B6",   x"7B",   x"EF",   x"22",   x"04",   x"C9",   x"5D",   x"90", 
  x"11",   x"DC",   x"48",   x"85",   x"A3",   x"6E",   x"FA",   x"37", 
  x"93",   x"5E",   x"CA",   x"07",   x"21",   x"EC",   x"78",   x"B5", 
  x"34",   x"F9",   x"6D",   x"A0",   x"86",   x"4B",   x"DF",   x"12", 
  x"1E",   x"D3",   x"47",   x"8A",   x"AC",   x"61",   x"F5",   x"38", 
  x"B9",   x"74",   x"E0",   x"2D",   x"0B",   x"C6",   x"52",   x"9F", 
  x"4A",   x"87",   x"13",   x"DE",   x"F8",   x"35",   x"A1",   x"6C", 
  x"ED",   x"20",   x"B4",   x"79",   x"5F",   x"92",   x"06",   x"CB", 
  x"C7",   x"0A",   x"9E",   x"53",   x"75",   x"B8",   x"2C",   x"E1", 
  x"60",   x"AD",   x"39",   x"F4",   x"D2",   x"1F",   x"8B",   x"46", 
  x"00",   x"CE",   x"5F",   x"91",   x"BE",   x"70",   x"E1",   x"2F", 
  x"BF",   x"71",   x"E0",   x"2E",   x"01",   x"CF",   x"5E",   x"90", 
  x"BD",   x"73",   x"E2",   x"2C",   x"03",   x"CD",   x"5C",   x"92", 
  x"02",   x"CC",   x"5D",   x"93",   x"BC",   x"72",   x"E3",   x"2D", 
  x"B9",   x"77",   x"E6",   x"28",   x"07",   x"C9",   x"58",   x"96", 
  x"06",   x"C8",   x"59",   x"97",   x"B8",   x"76",   x"E7",   x"29", 
  x"04",   x"CA",   x"5B",   x"95",   x"BA",   x"74",   x"E5",   x"2B", 
  x"BB",   x"75",   x"E4",   x"2A",   x"05",   x"CB",   x"5A",   x"94", 
  x"B1",   x"7F",   x"EE",   x"20",   x"0F",   x"C1",   x"50",   x"9E", 
  x"0E",   x"C0",   x"51",   x"9F",   x"B0",   x"7E",   x"EF",   x"21", 
  x"0C",   x"C2",   x"53",   x"9D",   x"B2",   x"7C",   x"ED",   x"23", 
  x"B3",   x"7D",   x"EC",   x"22",   x"0D",   x"C3",   x"52",   x"9C", 
  x"08",   x"C6",   x"57",   x"99",   x"B6",   x"78",   x"E9",   x"27", 
  x"B7",   x"79",   x"E8",   x"26",   x"09",   x"C7",   x"56",   x"98", 
  x"B5",   x"7B",   x"EA",   x"24",   x"0B",   x"C5",   x"54",   x"9A", 
  x"0A",   x"C4",   x"55",   x"9B",   x"B4",   x"7A",   x"EB",   x"25", 
  x"A1",   x"6F",   x"FE",   x"30",   x"1F",   x"D1",   x"40",   x"8E", 
  x"1E",   x"D0",   x"41",   x"8F",   x"A0",   x"6E",   x"FF",   x"31", 
  x"1C",   x"D2",   x"43",   x"8D",   x"A2",   x"6C",   x"FD",   x"33", 
  x"A3",   x"6D",   x"FC",   x"32",   x"1D",   x"D3",   x"42",   x"8C", 
  x"18",   x"D6",   x"47",   x"89",   x"A6",   x"68",   x"F9",   x"37", 
  x"A7",   x"69",   x"F8",   x"36",   x"19",   x"D7",   x"46",   x"88", 
  x"A5",   x"6B",   x"FA",   x"34",   x"1B",   x"D5",   x"44",   x"8A", 
  x"1A",   x"D4",   x"45",   x"8B",   x"A4",   x"6A",   x"FB",   x"35", 
  x"10",   x"DE",   x"4F",   x"81",   x"AE",   x"60",   x"F1",   x"3F", 
  x"AF",   x"61",   x"F0",   x"3E",   x"11",   x"DF",   x"4E",   x"80", 
  x"AD",   x"63",   x"F2",   x"3C",   x"13",   x"DD",   x"4C",   x"82", 
  x"12",   x"DC",   x"4D",   x"83",   x"AC",   x"62",   x"F3",   x"3D", 
  x"A9",   x"67",   x"F6",   x"38",   x"17",   x"D9",   x"48",   x"86", 
  x"16",   x"D8",   x"49",   x"87",   x"A8",   x"66",   x"F7",   x"39", 
  x"14",   x"DA",   x"4B",   x"85",   x"AA",   x"64",   x"F5",   x"3B", 
  x"AB",   x"65",   x"F4",   x"3A",   x"15",   x"DB",   x"4A",   x"84", 
  x"00",   x"CF",   x"5D",   x"92",   x"BA",   x"75",   x"E7",   x"28", 
  x"B7",   x"78",   x"EA",   x"25",   x"0D",   x"C2",   x"50",   x"9F", 
  x"AD",   x"62",   x"F0",   x"3F",   x"17",   x"D8",   x"4A",   x"85", 
  x"1A",   x"D5",   x"47",   x"88",   x"A0",   x"6F",   x"FD",   x"32", 
  x"99",   x"56",   x"C4",   x"0B",   x"23",   x"EC",   x"7E",   x"B1", 
  x"2E",   x"E1",   x"73",   x"BC",   x"94",   x"5B",   x"C9",   x"06", 
  x"34",   x"FB",   x"69",   x"A6",   x"8E",   x"41",   x"D3",   x"1C", 
  x"83",   x"4C",   x"DE",   x"11",   x"39",   x"F6",   x"64",   x"AB", 
  x"F1",   x"3E",   x"AC",   x"63",   x"4B",   x"84",   x"16",   x"D9", 
  x"46",   x"89",   x"1B",   x"D4",   x"FC",   x"33",   x"A1",   x"6E", 
  x"5C",   x"93",   x"01",   x"CE",   x"E6",   x"29",   x"BB",   x"74", 
  x"EB",   x"24",   x"B6",   x"79",   x"51",   x"9E",   x"0C",   x"C3", 
  x"68",   x"A7",   x"35",   x"FA",   x"D2",   x"1D",   x"8F",   x"40", 
  x"DF",   x"10",   x"82",   x"4D",   x"65",   x"AA",   x"38",   x"F7", 
  x"C5",   x"0A",   x"98",   x"57",   x"7F",   x"B0",   x"22",   x"ED", 
  x"72",   x"BD",   x"2F",   x"E0",   x"C8",   x"07",   x"95",   x"5A", 
  x"21",   x"EE",   x"7C",   x"B3",   x"9B",   x"54",   x"C6",   x"09", 
  x"96",   x"59",   x"CB",   x"04",   x"2C",   x"E3",   x"71",   x"BE", 
  x"8C",   x"43",   x"D1",   x"1E",   x"36",   x"F9",   x"6B",   x"A4", 
  x"3B",   x"F4",   x"66",   x"A9",   x"81",   x"4E",   x"DC",   x"13", 
  x"B8",   x"77",   x"E5",   x"2A",   x"02",   x"CD",   x"5F",   x"90", 
  x"0F",   x"C0",   x"52",   x"9D",   x"B5",   x"7A",   x"E8",   x"27", 
  x"15",   x"DA",   x"48",   x"87",   x"AF",   x"60",   x"F2",   x"3D", 
  x"A2",   x"6D",   x"FF",   x"30",   x"18",   x"D7",   x"45",   x"8A", 
  x"D0",   x"1F",   x"8D",   x"42",   x"6A",   x"A5",   x"37",   x"F8", 
  x"67",   x"A8",   x"3A",   x"F5",   x"DD",   x"12",   x"80",   x"4F", 
  x"7D",   x"B2",   x"20",   x"EF",   x"C7",   x"08",   x"9A",   x"55", 
  x"CA",   x"05",   x"97",   x"58",   x"70",   x"BF",   x"2D",   x"E2", 
  x"49",   x"86",   x"14",   x"DB",   x"F3",   x"3C",   x"AE",   x"61", 
  x"FE",   x"31",   x"A3",   x"6C",   x"44",   x"8B",   x"19",   x"D6", 
  x"E4",   x"2B",   x"B9",   x"76",   x"5E",   x"91",   x"03",   x"CC", 
  x"53",   x"9C",   x"0E",   x"C1",   x"E9",   x"26",   x"B4",   x"7B", 
  x"00",   x"D0",   x"63",   x"B3",   x"C6",   x"16",   x"A5",   x"75", 
  x"4F",   x"9F",   x"2C",   x"FC",   x"89",   x"59",   x"EA",   x"3A", 
  x"9E",   x"4E",   x"FD",   x"2D",   x"58",   x"88",   x"3B",   x"EB", 
  x"D1",   x"01",   x"B2",   x"62",   x"17",   x"C7",   x"74",   x"A4", 
  x"FF",   x"2F",   x"9C",   x"4C",   x"39",   x"E9",   x"5A",   x"8A", 
  x"B0",   x"60",   x"D3",   x"03",   x"76",   x"A6",   x"15",   x"C5", 
  x"61",   x"B1",   x"02",   x"D2",   x"A7",   x"77",   x"C4",   x"14", 
  x"2E",   x"FE",   x"4D",   x"9D",   x"E8",   x"38",   x"8B",   x"5B", 
  x"3D",   x"ED",   x"5E",   x"8E",   x"FB",   x"2B",   x"98",   x"48", 
  x"72",   x"A2",   x"11",   x"C1",   x"B4",   x"64",   x"D7",   x"07", 
  x"A3",   x"73",   x"C0",   x"10",   x"65",   x"B5",   x"06",   x"D6", 
  x"EC",   x"3C",   x"8F",   x"5F",   x"2A",   x"FA",   x"49",   x"99", 
  x"C2",   x"12",   x"A1",   x"71",   x"04",   x"D4",   x"67",   x"B7", 
  x"8D",   x"5D",   x"EE",   x"3E",   x"4B",   x"9B",   x"28",   x"F8", 
  x"5C",   x"8C",   x"3F",   x"EF",   x"9A",   x"4A",   x"F9",   x"29", 
  x"13",   x"C3",   x"70",   x"A0",   x"D5",   x"05",   x"B6",   x"66", 
  x"7A",   x"AA",   x"19",   x"C9",   x"BC",   x"6C",   x"DF",   x"0F", 
  x"35",   x"E5",   x"56",   x"86",   x"F3",   x"23",   x"90",   x"40", 
  x"E4",   x"34",   x"87",   x"57",   x"22",   x"F2",   x"41",   x"91", 
  x"AB",   x"7B",   x"C8",   x"18",   x"6D",   x"BD",   x"0E",   x"DE", 
  x"85",   x"55",   x"E6",   x"36",   x"43",   x"93",   x"20",   x"F0", 
  x"CA",   x"1A",   x"A9",   x"79",   x"0C",   x"DC",   x"6F",   x"BF", 
  x"1B",   x"CB",   x"78",   x"A8",   x"DD",   x"0D",   x"BE",   x"6E", 
  x"54",   x"84",   x"37",   x"E7",   x"92",   x"42",   x"F1",   x"21", 
  x"47",   x"97",   x"24",   x"F4",   x"81",   x"51",   x"E2",   x"32", 
  x"08",   x"D8",   x"6B",   x"BB",   x"CE",   x"1E",   x"AD",   x"7D", 
  x"D9",   x"09",   x"BA",   x"6A",   x"1F",   x"CF",   x"7C",   x"AC", 
  x"96",   x"46",   x"F5",   x"25",   x"50",   x"80",   x"33",   x"E3", 
  x"B8",   x"68",   x"DB",   x"0B",   x"7E",   x"AE",   x"1D",   x"CD", 
  x"F7",   x"27",   x"94",   x"44",   x"31",   x"E1",   x"52",   x"82", 
  x"26",   x"F6",   x"45",   x"95",   x"E0",   x"30",   x"83",   x"53", 
  x"69",   x"B9",   x"0A",   x"DA",   x"AF",   x"7F",   x"CC",   x"1C", 
  x"00",   x"D1",   x"61",   x"B0",   x"C2",   x"13",   x"A3",   x"72", 
  x"47",   x"96",   x"26",   x"F7",   x"85",   x"54",   x"E4",   x"35", 
  x"8E",   x"5F",   x"EF",   x"3E",   x"4C",   x"9D",   x"2D",   x"FC", 
  x"C9",   x"18",   x"A8",   x"79",   x"0B",   x"DA",   x"6A",   x"BB", 
  x"DF",   x"0E",   x"BE",   x"6F",   x"1D",   x"CC",   x"7C",   x"AD", 
  x"98",   x"49",   x"F9",   x"28",   x"5A",   x"8B",   x"3B",   x"EA", 
  x"51",   x"80",   x"30",   x"E1",   x"93",   x"42",   x"F2",   x"23", 
  x"16",   x"C7",   x"77",   x"A6",   x"D4",   x"05",   x"B5",   x"64", 
  x"7D",   x"AC",   x"1C",   x"CD",   x"BF",   x"6E",   x"DE",   x"0F", 
  x"3A",   x"EB",   x"5B",   x"8A",   x"F8",   x"29",   x"99",   x"48", 
  x"F3",   x"22",   x"92",   x"43",   x"31",   x"E0",   x"50",   x"81", 
  x"B4",   x"65",   x"D5",   x"04",   x"76",   x"A7",   x"17",   x"C6", 
  x"A2",   x"73",   x"C3",   x"12",   x"60",   x"B1",   x"01",   x"D0", 
  x"E5",   x"34",   x"84",   x"55",   x"27",   x"F6",   x"46",   x"97", 
  x"2C",   x"FD",   x"4D",   x"9C",   x"EE",   x"3F",   x"8F",   x"5E", 
  x"6B",   x"BA",   x"0A",   x"DB",   x"A9",   x"78",   x"C8",   x"19", 
  x"FA",   x"2B",   x"9B",   x"4A",   x"38",   x"E9",   x"59",   x"88", 
  x"BD",   x"6C",   x"DC",   x"0D",   x"7F",   x"AE",   x"1E",   x"CF", 
  x"74",   x"A5",   x"15",   x"C4",   x"B6",   x"67",   x"D7",   x"06", 
  x"33",   x"E2",   x"52",   x"83",   x"F1",   x"20",   x"90",   x"41", 
  x"25",   x"F4",   x"44",   x"95",   x"E7",   x"36",   x"86",   x"57", 
  x"62",   x"B3",   x"03",   x"D2",   x"A0",   x"71",   x"C1",   x"10", 
  x"AB",   x"7A",   x"CA",   x"1B",   x"69",   x"B8",   x"08",   x"D9", 
  x"EC",   x"3D",   x"8D",   x"5C",   x"2E",   x"FF",   x"4F",   x"9E", 
  x"87",   x"56",   x"E6",   x"37",   x"45",   x"94",   x"24",   x"F5", 
  x"C0",   x"11",   x"A1",   x"70",   x"02",   x"D3",   x"63",   x"B2", 
  x"09",   x"D8",   x"68",   x"B9",   x"CB",   x"1A",   x"AA",   x"7B", 
  x"4E",   x"9F",   x"2F",   x"FE",   x"8C",   x"5D",   x"ED",   x"3C", 
  x"58",   x"89",   x"39",   x"E8",   x"9A",   x"4B",   x"FB",   x"2A", 
  x"1F",   x"CE",   x"7E",   x"AF",   x"DD",   x"0C",   x"BC",   x"6D", 
  x"D6",   x"07",   x"B7",   x"66",   x"14",   x"C5",   x"75",   x"A4", 
  x"91",   x"40",   x"F0",   x"21",   x"53",   x"82",   x"32",   x"E3", 
  x"00",   x"D2",   x"67",   x"B5",   x"CE",   x"1C",   x"A9",   x"7B", 
  x"5F",   x"8D",   x"38",   x"EA",   x"91",   x"43",   x"F6",   x"24", 
  x"BE",   x"6C",   x"D9",   x"0B",   x"70",   x"A2",   x"17",   x"C5", 
  x"E1",   x"33",   x"86",   x"54",   x"2F",   x"FD",   x"48",   x"9A", 
  x"BF",   x"6D",   x"D8",   x"0A",   x"71",   x"A3",   x"16",   x"C4", 
  x"E0",   x"32",   x"87",   x"55",   x"2E",   x"FC",   x"49",   x"9B", 
  x"01",   x"D3",   x"66",   x"B4",   x"CF",   x"1D",   x"A8",   x"7A", 
  x"5E",   x"8C",   x"39",   x"EB",   x"90",   x"42",   x"F7",   x"25", 
  x"BD",   x"6F",   x"DA",   x"08",   x"73",   x"A1",   x"14",   x"C6", 
  x"E2",   x"30",   x"85",   x"57",   x"2C",   x"FE",   x"4B",   x"99", 
  x"03",   x"D1",   x"64",   x"B6",   x"CD",   x"1F",   x"AA",   x"78", 
  x"5C",   x"8E",   x"3B",   x"E9",   x"92",   x"40",   x"F5",   x"27", 
  x"02",   x"D0",   x"65",   x"B7",   x"CC",   x"1E",   x"AB",   x"79", 
  x"5D",   x"8F",   x"3A",   x"E8",   x"93",   x"41",   x"F4",   x"26", 
  x"BC",   x"6E",   x"DB",   x"09",   x"72",   x"A0",   x"15",   x"C7", 
  x"E3",   x"31",   x"84",   x"56",   x"2D",   x"FF",   x"4A",   x"98", 
  x"B9",   x"6B",   x"DE",   x"0C",   x"77",   x"A5",   x"10",   x"C2", 
  x"E6",   x"34",   x"81",   x"53",   x"28",   x"FA",   x"4F",   x"9D", 
  x"07",   x"D5",   x"60",   x"B2",   x"C9",   x"1B",   x"AE",   x"7C", 
  x"58",   x"8A",   x"3F",   x"ED",   x"96",   x"44",   x"F1",   x"23", 
  x"06",   x"D4",   x"61",   x"B3",   x"C8",   x"1A",   x"AF",   x"7D", 
  x"59",   x"8B",   x"3E",   x"EC",   x"97",   x"45",   x"F0",   x"22", 
  x"B8",   x"6A",   x"DF",   x"0D",   x"76",   x"A4",   x"11",   x"C3", 
  x"E7",   x"35",   x"80",   x"52",   x"29",   x"FB",   x"4E",   x"9C", 
  x"04",   x"D6",   x"63",   x"B1",   x"CA",   x"18",   x"AD",   x"7F", 
  x"5B",   x"89",   x"3C",   x"EE",   x"95",   x"47",   x"F2",   x"20", 
  x"BA",   x"68",   x"DD",   x"0F",   x"74",   x"A6",   x"13",   x"C1", 
  x"E5",   x"37",   x"82",   x"50",   x"2B",   x"F9",   x"4C",   x"9E", 
  x"BB",   x"69",   x"DC",   x"0E",   x"75",   x"A7",   x"12",   x"C0", 
  x"E4",   x"36",   x"83",   x"51",   x"2A",   x"F8",   x"4D",   x"9F", 
  x"05",   x"D7",   x"62",   x"B0",   x"CB",   x"19",   x"AC",   x"7E", 
  x"5A",   x"88",   x"3D",   x"EF",   x"94",   x"46",   x"F3",   x"21", 
  x"00",   x"D3",   x"65",   x"B6",   x"CA",   x"19",   x"AF",   x"7C", 
  x"57",   x"84",   x"32",   x"E1",   x"9D",   x"4E",   x"F8",   x"2B", 
  x"AE",   x"7D",   x"CB",   x"18",   x"64",   x"B7",   x"01",   x"D2", 
  x"F9",   x"2A",   x"9C",   x"4F",   x"33",   x"E0",   x"56",   x"85", 
  x"9F",   x"4C",   x"FA",   x"29",   x"55",   x"86",   x"30",   x"E3", 
  x"C8",   x"1B",   x"AD",   x"7E",   x"02",   x"D1",   x"67",   x"B4", 
  x"31",   x"E2",   x"54",   x"87",   x"FB",   x"28",   x"9E",   x"4D", 
  x"66",   x"B5",   x"03",   x"D0",   x"AC",   x"7F",   x"C9",   x"1A", 
  x"FD",   x"2E",   x"98",   x"4B",   x"37",   x"E4",   x"52",   x"81", 
  x"AA",   x"79",   x"CF",   x"1C",   x"60",   x"B3",   x"05",   x"D6", 
  x"53",   x"80",   x"36",   x"E5",   x"99",   x"4A",   x"FC",   x"2F", 
  x"04",   x"D7",   x"61",   x"B2",   x"CE",   x"1D",   x"AB",   x"78", 
  x"62",   x"B1",   x"07",   x"D4",   x"A8",   x"7B",   x"CD",   x"1E", 
  x"35",   x"E6",   x"50",   x"83",   x"FF",   x"2C",   x"9A",   x"49", 
  x"CC",   x"1F",   x"A9",   x"7A",   x"06",   x"D5",   x"63",   x"B0", 
  x"9B",   x"48",   x"FE",   x"2D",   x"51",   x"82",   x"34",   x"E7", 
  x"39",   x"EA",   x"5C",   x"8F",   x"F3",   x"20",   x"96",   x"45", 
  x"6E",   x"BD",   x"0B",   x"D8",   x"A4",   x"77",   x"C1",   x"12", 
  x"97",   x"44",   x"F2",   x"21",   x"5D",   x"8E",   x"38",   x"EB", 
  x"C0",   x"13",   x"A5",   x"76",   x"0A",   x"D9",   x"6F",   x"BC", 
  x"A6",   x"75",   x"C3",   x"10",   x"6C",   x"BF",   x"09",   x"DA", 
  x"F1",   x"22",   x"94",   x"47",   x"3B",   x"E8",   x"5E",   x"8D", 
  x"08",   x"DB",   x"6D",   x"BE",   x"C2",   x"11",   x"A7",   x"74", 
  x"5F",   x"8C",   x"3A",   x"E9",   x"95",   x"46",   x"F0",   x"23", 
  x"C4",   x"17",   x"A1",   x"72",   x"0E",   x"DD",   x"6B",   x"B8", 
  x"93",   x"40",   x"F6",   x"25",   x"59",   x"8A",   x"3C",   x"EF", 
  x"6A",   x"B9",   x"0F",   x"DC",   x"A0",   x"73",   x"C5",   x"16", 
  x"3D",   x"EE",   x"58",   x"8B",   x"F7",   x"24",   x"92",   x"41", 
  x"5B",   x"88",   x"3E",   x"ED",   x"91",   x"42",   x"F4",   x"27", 
  x"0C",   x"DF",   x"69",   x"BA",   x"C6",   x"15",   x"A3",   x"70", 
  x"F5",   x"26",   x"90",   x"43",   x"3F",   x"EC",   x"5A",   x"89", 
  x"A2",   x"71",   x"C7",   x"14",   x"68",   x"BB",   x"0D",   x"DE", 
  x"00",   x"D4",   x"6B",   x"BF",   x"D6",   x"02",   x"BD",   x"69", 
  x"6F",   x"BB",   x"04",   x"D0",   x"B9",   x"6D",   x"D2",   x"06", 
  x"DE",   x"0A",   x"B5",   x"61",   x"08",   x"DC",   x"63",   x"B7", 
  x"B1",   x"65",   x"DA",   x"0E",   x"67",   x"B3",   x"0C",   x"D8", 
  x"7F",   x"AB",   x"14",   x"C0",   x"A9",   x"7D",   x"C2",   x"16", 
  x"10",   x"C4",   x"7B",   x"AF",   x"C6",   x"12",   x"AD",   x"79", 
  x"A1",   x"75",   x"CA",   x"1E",   x"77",   x"A3",   x"1C",   x"C8", 
  x"CE",   x"1A",   x"A5",   x"71",   x"18",   x"CC",   x"73",   x"A7", 
  x"FE",   x"2A",   x"95",   x"41",   x"28",   x"FC",   x"43",   x"97", 
  x"91",   x"45",   x"FA",   x"2E",   x"47",   x"93",   x"2C",   x"F8", 
  x"20",   x"F4",   x"4B",   x"9F",   x"F6",   x"22",   x"9D",   x"49", 
  x"4F",   x"9B",   x"24",   x"F0",   x"99",   x"4D",   x"F2",   x"26", 
  x"81",   x"55",   x"EA",   x"3E",   x"57",   x"83",   x"3C",   x"E8", 
  x"EE",   x"3A",   x"85",   x"51",   x"38",   x"EC",   x"53",   x"87", 
  x"5F",   x"8B",   x"34",   x"E0",   x"89",   x"5D",   x"E2",   x"36", 
  x"30",   x"E4",   x"5B",   x"8F",   x"E6",   x"32",   x"8D",   x"59", 
  x"3F",   x"EB",   x"54",   x"80",   x"E9",   x"3D",   x"82",   x"56", 
  x"50",   x"84",   x"3B",   x"EF",   x"86",   x"52",   x"ED",   x"39", 
  x"E1",   x"35",   x"8A",   x"5E",   x"37",   x"E3",   x"5C",   x"88", 
  x"8E",   x"5A",   x"E5",   x"31",   x"58",   x"8C",   x"33",   x"E7", 
  x"40",   x"94",   x"2B",   x"FF",   x"96",   x"42",   x"FD",   x"29", 
  x"2F",   x"FB",   x"44",   x"90",   x"F9",   x"2D",   x"92",   x"46", 
  x"9E",   x"4A",   x"F5",   x"21",   x"48",   x"9C",   x"23",   x"F7", 
  x"F1",   x"25",   x"9A",   x"4E",   x"27",   x"F3",   x"4C",   x"98", 
  x"C1",   x"15",   x"AA",   x"7E",   x"17",   x"C3",   x"7C",   x"A8", 
  x"AE",   x"7A",   x"C5",   x"11",   x"78",   x"AC",   x"13",   x"C7", 
  x"1F",   x"CB",   x"74",   x"A0",   x"C9",   x"1D",   x"A2",   x"76", 
  x"70",   x"A4",   x"1B",   x"CF",   x"A6",   x"72",   x"CD",   x"19", 
  x"BE",   x"6A",   x"D5",   x"01",   x"68",   x"BC",   x"03",   x"D7", 
  x"D1",   x"05",   x"BA",   x"6E",   x"07",   x"D3",   x"6C",   x"B8", 
  x"60",   x"B4",   x"0B",   x"DF",   x"B6",   x"62",   x"DD",   x"09", 
  x"0F",   x"DB",   x"64",   x"B0",   x"D9",   x"0D",   x"B2",   x"66", 
  x"00",   x"D5",   x"69",   x"BC",   x"D2",   x"07",   x"BB",   x"6E", 
  x"67",   x"B2",   x"0E",   x"DB",   x"B5",   x"60",   x"DC",   x"09", 
  x"CE",   x"1B",   x"A7",   x"72",   x"1C",   x"C9",   x"75",   x"A0", 
  x"A9",   x"7C",   x"C0",   x"15",   x"7B",   x"AE",   x"12",   x"C7", 
  x"5F",   x"8A",   x"36",   x"E3",   x"8D",   x"58",   x"E4",   x"31", 
  x"38",   x"ED",   x"51",   x"84",   x"EA",   x"3F",   x"83",   x"56", 
  x"91",   x"44",   x"F8",   x"2D",   x"43",   x"96",   x"2A",   x"FF", 
  x"F6",   x"23",   x"9F",   x"4A",   x"24",   x"F1",   x"4D",   x"98", 
  x"BE",   x"6B",   x"D7",   x"02",   x"6C",   x"B9",   x"05",   x"D0", 
  x"D9",   x"0C",   x"B0",   x"65",   x"0B",   x"DE",   x"62",   x"B7", 
  x"70",   x"A5",   x"19",   x"CC",   x"A2",   x"77",   x"CB",   x"1E", 
  x"17",   x"C2",   x"7E",   x"AB",   x"C5",   x"10",   x"AC",   x"79", 
  x"E1",   x"34",   x"88",   x"5D",   x"33",   x"E6",   x"5A",   x"8F", 
  x"86",   x"53",   x"EF",   x"3A",   x"54",   x"81",   x"3D",   x"E8", 
  x"2F",   x"FA",   x"46",   x"93",   x"FD",   x"28",   x"94",   x"41", 
  x"48",   x"9D",   x"21",   x"F4",   x"9A",   x"4F",   x"F3",   x"26", 
  x"BF",   x"6A",   x"D6",   x"03",   x"6D",   x"B8",   x"04",   x"D1", 
  x"D8",   x"0D",   x"B1",   x"64",   x"0A",   x"DF",   x"63",   x"B6", 
  x"71",   x"A4",   x"18",   x"CD",   x"A3",   x"76",   x"CA",   x"1F", 
  x"16",   x"C3",   x"7F",   x"AA",   x"C4",   x"11",   x"AD",   x"78", 
  x"E0",   x"35",   x"89",   x"5C",   x"32",   x"E7",   x"5B",   x"8E", 
  x"87",   x"52",   x"EE",   x"3B",   x"55",   x"80",   x"3C",   x"E9", 
  x"2E",   x"FB",   x"47",   x"92",   x"FC",   x"29",   x"95",   x"40", 
  x"49",   x"9C",   x"20",   x"F5",   x"9B",   x"4E",   x"F2",   x"27", 
  x"01",   x"D4",   x"68",   x"BD",   x"D3",   x"06",   x"BA",   x"6F", 
  x"66",   x"B3",   x"0F",   x"DA",   x"B4",   x"61",   x"DD",   x"08", 
  x"CF",   x"1A",   x"A6",   x"73",   x"1D",   x"C8",   x"74",   x"A1", 
  x"A8",   x"7D",   x"C1",   x"14",   x"7A",   x"AF",   x"13",   x"C6", 
  x"5E",   x"8B",   x"37",   x"E2",   x"8C",   x"59",   x"E5",   x"30", 
  x"39",   x"EC",   x"50",   x"85",   x"EB",   x"3E",   x"82",   x"57", 
  x"90",   x"45",   x"F9",   x"2C",   x"42",   x"97",   x"2B",   x"FE", 
  x"F7",   x"22",   x"9E",   x"4B",   x"25",   x"F0",   x"4C",   x"99", 
  x"00",   x"D6",   x"6F",   x"B9",   x"DE",   x"08",   x"B1",   x"67", 
  x"7F",   x"A9",   x"10",   x"C6",   x"A1",   x"77",   x"CE",   x"18", 
  x"FE",   x"28",   x"91",   x"47",   x"20",   x"F6",   x"4F",   x"99", 
  x"81",   x"57",   x"EE",   x"38",   x"5F",   x"89",   x"30",   x"E6", 
  x"3F",   x"E9",   x"50",   x"86",   x"E1",   x"37",   x"8E",   x"58", 
  x"40",   x"96",   x"2F",   x"F9",   x"9E",   x"48",   x"F1",   x"27", 
  x"C1",   x"17",   x"AE",   x"78",   x"1F",   x"C9",   x"70",   x"A6", 
  x"BE",   x"68",   x"D1",   x"07",   x"60",   x"B6",   x"0F",   x"D9", 
  x"7E",   x"A8",   x"11",   x"C7",   x"A0",   x"76",   x"CF",   x"19", 
  x"01",   x"D7",   x"6E",   x"B8",   x"DF",   x"09",   x"B0",   x"66", 
  x"80",   x"56",   x"EF",   x"39",   x"5E",   x"88",   x"31",   x"E7", 
  x"FF",   x"29",   x"90",   x"46",   x"21",   x"F7",   x"4E",   x"98", 
  x"41",   x"97",   x"2E",   x"F8",   x"9F",   x"49",   x"F0",   x"26", 
  x"3E",   x"E8",   x"51",   x"87",   x"E0",   x"36",   x"8F",   x"59", 
  x"BF",   x"69",   x"D0",   x"06",   x"61",   x"B7",   x"0E",   x"D8", 
  x"C0",   x"16",   x"AF",   x"79",   x"1E",   x"C8",   x"71",   x"A7", 
  x"FC",   x"2A",   x"93",   x"45",   x"22",   x"F4",   x"4D",   x"9B", 
  x"83",   x"55",   x"EC",   x"3A",   x"5D",   x"8B",   x"32",   x"E4", 
  x"02",   x"D4",   x"6D",   x"BB",   x"DC",   x"0A",   x"B3",   x"65", 
  x"7D",   x"AB",   x"12",   x"C4",   x"A3",   x"75",   x"CC",   x"1A", 
  x"C3",   x"15",   x"AC",   x"7A",   x"1D",   x"CB",   x"72",   x"A4", 
  x"BC",   x"6A",   x"D3",   x"05",   x"62",   x"B4",   x"0D",   x"DB", 
  x"3D",   x"EB",   x"52",   x"84",   x"E3",   x"35",   x"8C",   x"5A", 
  x"42",   x"94",   x"2D",   x"FB",   x"9C",   x"4A",   x"F3",   x"25", 
  x"82",   x"54",   x"ED",   x"3B",   x"5C",   x"8A",   x"33",   x"E5", 
  x"FD",   x"2B",   x"92",   x"44",   x"23",   x"F5",   x"4C",   x"9A", 
  x"7C",   x"AA",   x"13",   x"C5",   x"A2",   x"74",   x"CD",   x"1B", 
  x"03",   x"D5",   x"6C",   x"BA",   x"DD",   x"0B",   x"B2",   x"64", 
  x"BD",   x"6B",   x"D2",   x"04",   x"63",   x"B5",   x"0C",   x"DA", 
  x"C2",   x"14",   x"AD",   x"7B",   x"1C",   x"CA",   x"73",   x"A5", 
  x"43",   x"95",   x"2C",   x"FA",   x"9D",   x"4B",   x"F2",   x"24", 
  x"3C",   x"EA",   x"53",   x"85",   x"E2",   x"34",   x"8D",   x"5B", 
  x"00",   x"D7",   x"6D",   x"BA",   x"DA",   x"0D",   x"B7",   x"60", 
  x"77",   x"A0",   x"1A",   x"CD",   x"AD",   x"7A",   x"C0",   x"17", 
  x"EE",   x"39",   x"83",   x"54",   x"34",   x"E3",   x"59",   x"8E", 
  x"99",   x"4E",   x"F4",   x"23",   x"43",   x"94",   x"2E",   x"F9", 
  x"1F",   x"C8",   x"72",   x"A5",   x"C5",   x"12",   x"A8",   x"7F", 
  x"68",   x"BF",   x"05",   x"D2",   x"B2",   x"65",   x"DF",   x"08", 
  x"F1",   x"26",   x"9C",   x"4B",   x"2B",   x"FC",   x"46",   x"91", 
  x"86",   x"51",   x"EB",   x"3C",   x"5C",   x"8B",   x"31",   x"E6", 
  x"3E",   x"E9",   x"53",   x"84",   x"E4",   x"33",   x"89",   x"5E", 
  x"49",   x"9E",   x"24",   x"F3",   x"93",   x"44",   x"FE",   x"29", 
  x"D0",   x"07",   x"BD",   x"6A",   x"0A",   x"DD",   x"67",   x"B0", 
  x"A7",   x"70",   x"CA",   x"1D",   x"7D",   x"AA",   x"10",   x"C7", 
  x"21",   x"F6",   x"4C",   x"9B",   x"FB",   x"2C",   x"96",   x"41", 
  x"56",   x"81",   x"3B",   x"EC",   x"8C",   x"5B",   x"E1",   x"36", 
  x"CF",   x"18",   x"A2",   x"75",   x"15",   x"C2",   x"78",   x"AF", 
  x"B8",   x"6F",   x"D5",   x"02",   x"62",   x"B5",   x"0F",   x"D8", 
  x"7C",   x"AB",   x"11",   x"C6",   x"A6",   x"71",   x"CB",   x"1C", 
  x"0B",   x"DC",   x"66",   x"B1",   x"D1",   x"06",   x"BC",   x"6B", 
  x"92",   x"45",   x"FF",   x"28",   x"48",   x"9F",   x"25",   x"F2", 
  x"E5",   x"32",   x"88",   x"5F",   x"3F",   x"E8",   x"52",   x"85", 
  x"63",   x"B4",   x"0E",   x"D9",   x"B9",   x"6E",   x"D4",   x"03", 
  x"14",   x"C3",   x"79",   x"AE",   x"CE",   x"19",   x"A3",   x"74", 
  x"8D",   x"5A",   x"E0",   x"37",   x"57",   x"80",   x"3A",   x"ED", 
  x"FA",   x"2D",   x"97",   x"40",   x"20",   x"F7",   x"4D",   x"9A", 
  x"42",   x"95",   x"2F",   x"F8",   x"98",   x"4F",   x"F5",   x"22", 
  x"35",   x"E2",   x"58",   x"8F",   x"EF",   x"38",   x"82",   x"55", 
  x"AC",   x"7B",   x"C1",   x"16",   x"76",   x"A1",   x"1B",   x"CC", 
  x"DB",   x"0C",   x"B6",   x"61",   x"01",   x"D6",   x"6C",   x"BB", 
  x"5D",   x"8A",   x"30",   x"E7",   x"87",   x"50",   x"EA",   x"3D", 
  x"2A",   x"FD",   x"47",   x"90",   x"F0",   x"27",   x"9D",   x"4A", 
  x"B3",   x"64",   x"DE",   x"09",   x"69",   x"BE",   x"04",   x"D3", 
  x"C4",   x"13",   x"A9",   x"7E",   x"1E",   x"C9",   x"73",   x"A4", 
  x"00",   x"D8",   x"73",   x"AB",   x"E6",   x"3E",   x"95",   x"4D", 
  x"0F",   x"D7",   x"7C",   x"A4",   x"E9",   x"31",   x"9A",   x"42", 
  x"1E",   x"C6",   x"6D",   x"B5",   x"F8",   x"20",   x"8B",   x"53", 
  x"11",   x"C9",   x"62",   x"BA",   x"F7",   x"2F",   x"84",   x"5C", 
  x"3C",   x"E4",   x"4F",   x"97",   x"DA",   x"02",   x"A9",   x"71", 
  x"33",   x"EB",   x"40",   x"98",   x"D5",   x"0D",   x"A6",   x"7E", 
  x"22",   x"FA",   x"51",   x"89",   x"C4",   x"1C",   x"B7",   x"6F", 
  x"2D",   x"F5",   x"5E",   x"86",   x"CB",   x"13",   x"B8",   x"60", 
  x"78",   x"A0",   x"0B",   x"D3",   x"9E",   x"46",   x"ED",   x"35", 
  x"77",   x"AF",   x"04",   x"DC",   x"91",   x"49",   x"E2",   x"3A", 
  x"66",   x"BE",   x"15",   x"CD",   x"80",   x"58",   x"F3",   x"2B", 
  x"69",   x"B1",   x"1A",   x"C2",   x"8F",   x"57",   x"FC",   x"24", 
  x"44",   x"9C",   x"37",   x"EF",   x"A2",   x"7A",   x"D1",   x"09", 
  x"4B",   x"93",   x"38",   x"E0",   x"AD",   x"75",   x"DE",   x"06", 
  x"5A",   x"82",   x"29",   x"F1",   x"BC",   x"64",   x"CF",   x"17", 
  x"55",   x"8D",   x"26",   x"FE",   x"B3",   x"6B",   x"C0",   x"18", 
  x"F0",   x"28",   x"83",   x"5B",   x"16",   x"CE",   x"65",   x"BD", 
  x"FF",   x"27",   x"8C",   x"54",   x"19",   x"C1",   x"6A",   x"B2", 
  x"EE",   x"36",   x"9D",   x"45",   x"08",   x"D0",   x"7B",   x"A3", 
  x"E1",   x"39",   x"92",   x"4A",   x"07",   x"DF",   x"74",   x"AC", 
  x"CC",   x"14",   x"BF",   x"67",   x"2A",   x"F2",   x"59",   x"81", 
  x"C3",   x"1B",   x"B0",   x"68",   x"25",   x"FD",   x"56",   x"8E", 
  x"D2",   x"0A",   x"A1",   x"79",   x"34",   x"EC",   x"47",   x"9F", 
  x"DD",   x"05",   x"AE",   x"76",   x"3B",   x"E3",   x"48",   x"90", 
  x"88",   x"50",   x"FB",   x"23",   x"6E",   x"B6",   x"1D",   x"C5", 
  x"87",   x"5F",   x"F4",   x"2C",   x"61",   x"B9",   x"12",   x"CA", 
  x"96",   x"4E",   x"E5",   x"3D",   x"70",   x"A8",   x"03",   x"DB", 
  x"99",   x"41",   x"EA",   x"32",   x"7F",   x"A7",   x"0C",   x"D4", 
  x"B4",   x"6C",   x"C7",   x"1F",   x"52",   x"8A",   x"21",   x"F9", 
  x"BB",   x"63",   x"C8",   x"10",   x"5D",   x"85",   x"2E",   x"F6", 
  x"AA",   x"72",   x"D9",   x"01",   x"4C",   x"94",   x"3F",   x"E7", 
  x"A5",   x"7D",   x"D6",   x"0E",   x"43",   x"9B",   x"30",   x"E8", 
  x"00",   x"D9",   x"71",   x"A8",   x"E2",   x"3B",   x"93",   x"4A", 
  x"07",   x"DE",   x"76",   x"AF",   x"E5",   x"3C",   x"94",   x"4D", 
  x"0E",   x"D7",   x"7F",   x"A6",   x"EC",   x"35",   x"9D",   x"44", 
  x"09",   x"D0",   x"78",   x"A1",   x"EB",   x"32",   x"9A",   x"43", 
  x"1C",   x"C5",   x"6D",   x"B4",   x"FE",   x"27",   x"8F",   x"56", 
  x"1B",   x"C2",   x"6A",   x"B3",   x"F9",   x"20",   x"88",   x"51", 
  x"12",   x"CB",   x"63",   x"BA",   x"F0",   x"29",   x"81",   x"58", 
  x"15",   x"CC",   x"64",   x"BD",   x"F7",   x"2E",   x"86",   x"5F", 
  x"38",   x"E1",   x"49",   x"90",   x"DA",   x"03",   x"AB",   x"72", 
  x"3F",   x"E6",   x"4E",   x"97",   x"DD",   x"04",   x"AC",   x"75", 
  x"36",   x"EF",   x"47",   x"9E",   x"D4",   x"0D",   x"A5",   x"7C", 
  x"31",   x"E8",   x"40",   x"99",   x"D3",   x"0A",   x"A2",   x"7B", 
  x"24",   x"FD",   x"55",   x"8C",   x"C6",   x"1F",   x"B7",   x"6E", 
  x"23",   x"FA",   x"52",   x"8B",   x"C1",   x"18",   x"B0",   x"69", 
  x"2A",   x"F3",   x"5B",   x"82",   x"C8",   x"11",   x"B9",   x"60", 
  x"2D",   x"F4",   x"5C",   x"85",   x"CF",   x"16",   x"BE",   x"67", 
  x"70",   x"A9",   x"01",   x"D8",   x"92",   x"4B",   x"E3",   x"3A", 
  x"77",   x"AE",   x"06",   x"DF",   x"95",   x"4C",   x"E4",   x"3D", 
  x"7E",   x"A7",   x"0F",   x"D6",   x"9C",   x"45",   x"ED",   x"34", 
  x"79",   x"A0",   x"08",   x"D1",   x"9B",   x"42",   x"EA",   x"33", 
  x"6C",   x"B5",   x"1D",   x"C4",   x"8E",   x"57",   x"FF",   x"26", 
  x"6B",   x"B2",   x"1A",   x"C3",   x"89",   x"50",   x"F8",   x"21", 
  x"62",   x"BB",   x"13",   x"CA",   x"80",   x"59",   x"F1",   x"28", 
  x"65",   x"BC",   x"14",   x"CD",   x"87",   x"5E",   x"F6",   x"2F", 
  x"48",   x"91",   x"39",   x"E0",   x"AA",   x"73",   x"DB",   x"02", 
  x"4F",   x"96",   x"3E",   x"E7",   x"AD",   x"74",   x"DC",   x"05", 
  x"46",   x"9F",   x"37",   x"EE",   x"A4",   x"7D",   x"D5",   x"0C", 
  x"41",   x"98",   x"30",   x"E9",   x"A3",   x"7A",   x"D2",   x"0B", 
  x"54",   x"8D",   x"25",   x"FC",   x"B6",   x"6F",   x"C7",   x"1E", 
  x"53",   x"8A",   x"22",   x"FB",   x"B1",   x"68",   x"C0",   x"19", 
  x"5A",   x"83",   x"2B",   x"F2",   x"B8",   x"61",   x"C9",   x"10", 
  x"5D",   x"84",   x"2C",   x"F5",   x"BF",   x"66",   x"CE",   x"17", 
  x"00",   x"DA",   x"77",   x"AD",   x"EE",   x"34",   x"99",   x"43", 
  x"1F",   x"C5",   x"68",   x"B2",   x"F1",   x"2B",   x"86",   x"5C", 
  x"3E",   x"E4",   x"49",   x"93",   x"D0",   x"0A",   x"A7",   x"7D", 
  x"21",   x"FB",   x"56",   x"8C",   x"CF",   x"15",   x"B8",   x"62", 
  x"7C",   x"A6",   x"0B",   x"D1",   x"92",   x"48",   x"E5",   x"3F", 
  x"63",   x"B9",   x"14",   x"CE",   x"8D",   x"57",   x"FA",   x"20", 
  x"42",   x"98",   x"35",   x"EF",   x"AC",   x"76",   x"DB",   x"01", 
  x"5D",   x"87",   x"2A",   x"F0",   x"B3",   x"69",   x"C4",   x"1E", 
  x"F8",   x"22",   x"8F",   x"55",   x"16",   x"CC",   x"61",   x"BB", 
  x"E7",   x"3D",   x"90",   x"4A",   x"09",   x"D3",   x"7E",   x"A4", 
  x"C6",   x"1C",   x"B1",   x"6B",   x"28",   x"F2",   x"5F",   x"85", 
  x"D9",   x"03",   x"AE",   x"74",   x"37",   x"ED",   x"40",   x"9A", 
  x"84",   x"5E",   x"F3",   x"29",   x"6A",   x"B0",   x"1D",   x"C7", 
  x"9B",   x"41",   x"EC",   x"36",   x"75",   x"AF",   x"02",   x"D8", 
  x"BA",   x"60",   x"CD",   x"17",   x"54",   x"8E",   x"23",   x"F9", 
  x"A5",   x"7F",   x"D2",   x"08",   x"4B",   x"91",   x"3C",   x"E6", 
  x"33",   x"E9",   x"44",   x"9E",   x"DD",   x"07",   x"AA",   x"70", 
  x"2C",   x"F6",   x"5B",   x"81",   x"C2",   x"18",   x"B5",   x"6F", 
  x"0D",   x"D7",   x"7A",   x"A0",   x"E3",   x"39",   x"94",   x"4E", 
  x"12",   x"C8",   x"65",   x"BF",   x"FC",   x"26",   x"8B",   x"51", 
  x"4F",   x"95",   x"38",   x"E2",   x"A1",   x"7B",   x"D6",   x"0C", 
  x"50",   x"8A",   x"27",   x"FD",   x"BE",   x"64",   x"C9",   x"13", 
  x"71",   x"AB",   x"06",   x"DC",   x"9F",   x"45",   x"E8",   x"32", 
  x"6E",   x"B4",   x"19",   x"C3",   x"80",   x"5A",   x"F7",   x"2D", 
  x"CB",   x"11",   x"BC",   x"66",   x"25",   x"FF",   x"52",   x"88", 
  x"D4",   x"0E",   x"A3",   x"79",   x"3A",   x"E0",   x"4D",   x"97", 
  x"F5",   x"2F",   x"82",   x"58",   x"1B",   x"C1",   x"6C",   x"B6", 
  x"EA",   x"30",   x"9D",   x"47",   x"04",   x"DE",   x"73",   x"A9", 
  x"B7",   x"6D",   x"C0",   x"1A",   x"59",   x"83",   x"2E",   x"F4", 
  x"A8",   x"72",   x"DF",   x"05",   x"46",   x"9C",   x"31",   x"EB", 
  x"89",   x"53",   x"FE",   x"24",   x"67",   x"BD",   x"10",   x"CA", 
  x"96",   x"4C",   x"E1",   x"3B",   x"78",   x"A2",   x"0F",   x"D5", 
  x"00",   x"DB",   x"75",   x"AE",   x"EA",   x"31",   x"9F",   x"44", 
  x"17",   x"CC",   x"62",   x"B9",   x"FD",   x"26",   x"88",   x"53", 
  x"2E",   x"F5",   x"5B",   x"80",   x"C4",   x"1F",   x"B1",   x"6A", 
  x"39",   x"E2",   x"4C",   x"97",   x"D3",   x"08",   x"A6",   x"7D", 
  x"5C",   x"87",   x"29",   x"F2",   x"B6",   x"6D",   x"C3",   x"18", 
  x"4B",   x"90",   x"3E",   x"E5",   x"A1",   x"7A",   x"D4",   x"0F", 
  x"72",   x"A9",   x"07",   x"DC",   x"98",   x"43",   x"ED",   x"36", 
  x"65",   x"BE",   x"10",   x"CB",   x"8F",   x"54",   x"FA",   x"21", 
  x"B8",   x"63",   x"CD",   x"16",   x"52",   x"89",   x"27",   x"FC", 
  x"AF",   x"74",   x"DA",   x"01",   x"45",   x"9E",   x"30",   x"EB", 
  x"96",   x"4D",   x"E3",   x"38",   x"7C",   x"A7",   x"09",   x"D2", 
  x"81",   x"5A",   x"F4",   x"2F",   x"6B",   x"B0",   x"1E",   x"C5", 
  x"E4",   x"3F",   x"91",   x"4A",   x"0E",   x"D5",   x"7B",   x"A0", 
  x"F3",   x"28",   x"86",   x"5D",   x"19",   x"C2",   x"6C",   x"B7", 
  x"CA",   x"11",   x"BF",   x"64",   x"20",   x"FB",   x"55",   x"8E", 
  x"DD",   x"06",   x"A8",   x"73",   x"37",   x"EC",   x"42",   x"99", 
  x"B3",   x"68",   x"C6",   x"1D",   x"59",   x"82",   x"2C",   x"F7", 
  x"A4",   x"7F",   x"D1",   x"0A",   x"4E",   x"95",   x"3B",   x"E0", 
  x"9D",   x"46",   x"E8",   x"33",   x"77",   x"AC",   x"02",   x"D9", 
  x"8A",   x"51",   x"FF",   x"24",   x"60",   x"BB",   x"15",   x"CE", 
  x"EF",   x"34",   x"9A",   x"41",   x"05",   x"DE",   x"70",   x"AB", 
  x"F8",   x"23",   x"8D",   x"56",   x"12",   x"C9",   x"67",   x"BC", 
  x"C1",   x"1A",   x"B4",   x"6F",   x"2B",   x"F0",   x"5E",   x"85", 
  x"D6",   x"0D",   x"A3",   x"78",   x"3C",   x"E7",   x"49",   x"92", 
  x"0B",   x"D0",   x"7E",   x"A5",   x"E1",   x"3A",   x"94",   x"4F", 
  x"1C",   x"C7",   x"69",   x"B2",   x"F6",   x"2D",   x"83",   x"58", 
  x"25",   x"FE",   x"50",   x"8B",   x"CF",   x"14",   x"BA",   x"61", 
  x"32",   x"E9",   x"47",   x"9C",   x"D8",   x"03",   x"AD",   x"76", 
  x"57",   x"8C",   x"22",   x"F9",   x"BD",   x"66",   x"C8",   x"13", 
  x"40",   x"9B",   x"35",   x"EE",   x"AA",   x"71",   x"DF",   x"04", 
  x"79",   x"A2",   x"0C",   x"D7",   x"93",   x"48",   x"E6",   x"3D", 
  x"6E",   x"B5",   x"1B",   x"C0",   x"84",   x"5F",   x"F1",   x"2A", 
  x"00",   x"DC",   x"7B",   x"A7",   x"F6",   x"2A",   x"8D",   x"51", 
  x"2F",   x"F3",   x"54",   x"88",   x"D9",   x"05",   x"A2",   x"7E", 
  x"5E",   x"82",   x"25",   x"F9",   x"A8",   x"74",   x"D3",   x"0F", 
  x"71",   x"AD",   x"0A",   x"D6",   x"87",   x"5B",   x"FC",   x"20", 
  x"BC",   x"60",   x"C7",   x"1B",   x"4A",   x"96",   x"31",   x"ED", 
  x"93",   x"4F",   x"E8",   x"34",   x"65",   x"B9",   x"1E",   x"C2", 
  x"E2",   x"3E",   x"99",   x"45",   x"14",   x"C8",   x"6F",   x"B3", 
  x"CD",   x"11",   x"B6",   x"6A",   x"3B",   x"E7",   x"40",   x"9C", 
  x"BB",   x"67",   x"C0",   x"1C",   x"4D",   x"91",   x"36",   x"EA", 
  x"94",   x"48",   x"EF",   x"33",   x"62",   x"BE",   x"19",   x"C5", 
  x"E5",   x"39",   x"9E",   x"42",   x"13",   x"CF",   x"68",   x"B4", 
  x"CA",   x"16",   x"B1",   x"6D",   x"3C",   x"E0",   x"47",   x"9B", 
  x"07",   x"DB",   x"7C",   x"A0",   x"F1",   x"2D",   x"8A",   x"56", 
  x"28",   x"F4",   x"53",   x"8F",   x"DE",   x"02",   x"A5",   x"79", 
  x"59",   x"85",   x"22",   x"FE",   x"AF",   x"73",   x"D4",   x"08", 
  x"76",   x"AA",   x"0D",   x"D1",   x"80",   x"5C",   x"FB",   x"27", 
  x"B5",   x"69",   x"CE",   x"12",   x"43",   x"9F",   x"38",   x"E4", 
  x"9A",   x"46",   x"E1",   x"3D",   x"6C",   x"B0",   x"17",   x"CB", 
  x"EB",   x"37",   x"90",   x"4C",   x"1D",   x"C1",   x"66",   x"BA", 
  x"C4",   x"18",   x"BF",   x"63",   x"32",   x"EE",   x"49",   x"95", 
  x"09",   x"D5",   x"72",   x"AE",   x"FF",   x"23",   x"84",   x"58", 
  x"26",   x"FA",   x"5D",   x"81",   x"D0",   x"0C",   x"AB",   x"77", 
  x"57",   x"8B",   x"2C",   x"F0",   x"A1",   x"7D",   x"DA",   x"06", 
  x"78",   x"A4",   x"03",   x"DF",   x"8E",   x"52",   x"F5",   x"29", 
  x"0E",   x"D2",   x"75",   x"A9",   x"F8",   x"24",   x"83",   x"5F", 
  x"21",   x"FD",   x"5A",   x"86",   x"D7",   x"0B",   x"AC",   x"70", 
  x"50",   x"8C",   x"2B",   x"F7",   x"A6",   x"7A",   x"DD",   x"01", 
  x"7F",   x"A3",   x"04",   x"D8",   x"89",   x"55",   x"F2",   x"2E", 
  x"B2",   x"6E",   x"C9",   x"15",   x"44",   x"98",   x"3F",   x"E3", 
  x"9D",   x"41",   x"E6",   x"3A",   x"6B",   x"B7",   x"10",   x"CC", 
  x"EC",   x"30",   x"97",   x"4B",   x"1A",   x"C6",   x"61",   x"BD", 
  x"C3",   x"1F",   x"B8",   x"64",   x"35",   x"E9",   x"4E",   x"92", 
  x"00",   x"DD",   x"79",   x"A4",   x"F2",   x"2F",   x"8B",   x"56", 
  x"27",   x"FA",   x"5E",   x"83",   x"D5",   x"08",   x"AC",   x"71", 
  x"4E",   x"93",   x"37",   x"EA",   x"BC",   x"61",   x"C5",   x"18", 
  x"69",   x"B4",   x"10",   x"CD",   x"9B",   x"46",   x"E2",   x"3F", 
  x"9C",   x"41",   x"E5",   x"38",   x"6E",   x"B3",   x"17",   x"CA", 
  x"BB",   x"66",   x"C2",   x"1F",   x"49",   x"94",   x"30",   x"ED", 
  x"D2",   x"0F",   x"AB",   x"76",   x"20",   x"FD",   x"59",   x"84", 
  x"F5",   x"28",   x"8C",   x"51",   x"07",   x"DA",   x"7E",   x"A3", 
  x"FB",   x"26",   x"82",   x"5F",   x"09",   x"D4",   x"70",   x"AD", 
  x"DC",   x"01",   x"A5",   x"78",   x"2E",   x"F3",   x"57",   x"8A", 
  x"B5",   x"68",   x"CC",   x"11",   x"47",   x"9A",   x"3E",   x"E3", 
  x"92",   x"4F",   x"EB",   x"36",   x"60",   x"BD",   x"19",   x"C4", 
  x"67",   x"BA",   x"1E",   x"C3",   x"95",   x"48",   x"EC",   x"31", 
  x"40",   x"9D",   x"39",   x"E4",   x"B2",   x"6F",   x"CB",   x"16", 
  x"29",   x"F4",   x"50",   x"8D",   x"DB",   x"06",   x"A2",   x"7F", 
  x"0E",   x"D3",   x"77",   x"AA",   x"FC",   x"21",   x"85",   x"58", 
  x"35",   x"E8",   x"4C",   x"91",   x"C7",   x"1A",   x"BE",   x"63", 
  x"12",   x"CF",   x"6B",   x"B6",   x"E0",   x"3D",   x"99",   x"44", 
  x"7B",   x"A6",   x"02",   x"DF",   x"89",   x"54",   x"F0",   x"2D", 
  x"5C",   x"81",   x"25",   x"F8",   x"AE",   x"73",   x"D7",   x"0A", 
  x"A9",   x"74",   x"D0",   x"0D",   x"5B",   x"86",   x"22",   x"FF", 
  x"8E",   x"53",   x"F7",   x"2A",   x"7C",   x"A1",   x"05",   x"D8", 
  x"E7",   x"3A",   x"9E",   x"43",   x"15",   x"C8",   x"6C",   x"B1", 
  x"C0",   x"1D",   x"B9",   x"64",   x"32",   x"EF",   x"4B",   x"96", 
  x"CE",   x"13",   x"B7",   x"6A",   x"3C",   x"E1",   x"45",   x"98", 
  x"E9",   x"34",   x"90",   x"4D",   x"1B",   x"C6",   x"62",   x"BF", 
  x"80",   x"5D",   x"F9",   x"24",   x"72",   x"AF",   x"0B",   x"D6", 
  x"A7",   x"7A",   x"DE",   x"03",   x"55",   x"88",   x"2C",   x"F1", 
  x"52",   x"8F",   x"2B",   x"F6",   x"A0",   x"7D",   x"D9",   x"04", 
  x"75",   x"A8",   x"0C",   x"D1",   x"87",   x"5A",   x"FE",   x"23", 
  x"1C",   x"C1",   x"65",   x"B8",   x"EE",   x"33",   x"97",   x"4A", 
  x"3B",   x"E6",   x"42",   x"9F",   x"C9",   x"14",   x"B0",   x"6D", 
  x"00",   x"DE",   x"7F",   x"A1",   x"FE",   x"20",   x"81",   x"5F", 
  x"3F",   x"E1",   x"40",   x"9E",   x"C1",   x"1F",   x"BE",   x"60", 
  x"7E",   x"A0",   x"01",   x"DF",   x"80",   x"5E",   x"FF",   x"21", 
  x"41",   x"9F",   x"3E",   x"E0",   x"BF",   x"61",   x"C0",   x"1E", 
  x"FC",   x"22",   x"83",   x"5D",   x"02",   x"DC",   x"7D",   x"A3", 
  x"C3",   x"1D",   x"BC",   x"62",   x"3D",   x"E3",   x"42",   x"9C", 
  x"82",   x"5C",   x"FD",   x"23",   x"7C",   x"A2",   x"03",   x"DD", 
  x"BD",   x"63",   x"C2",   x"1C",   x"43",   x"9D",   x"3C",   x"E2", 
  x"3B",   x"E5",   x"44",   x"9A",   x"C5",   x"1B",   x"BA",   x"64", 
  x"04",   x"DA",   x"7B",   x"A5",   x"FA",   x"24",   x"85",   x"5B", 
  x"45",   x"9B",   x"3A",   x"E4",   x"BB",   x"65",   x"C4",   x"1A", 
  x"7A",   x"A4",   x"05",   x"DB",   x"84",   x"5A",   x"FB",   x"25", 
  x"C7",   x"19",   x"B8",   x"66",   x"39",   x"E7",   x"46",   x"98", 
  x"F8",   x"26",   x"87",   x"59",   x"06",   x"D8",   x"79",   x"A7", 
  x"B9",   x"67",   x"C6",   x"18",   x"47",   x"99",   x"38",   x"E6", 
  x"86",   x"58",   x"F9",   x"27",   x"78",   x"A6",   x"07",   x"D9", 
  x"76",   x"A8",   x"09",   x"D7",   x"88",   x"56",   x"F7",   x"29", 
  x"49",   x"97",   x"36",   x"E8",   x"B7",   x"69",   x"C8",   x"16", 
  x"08",   x"D6",   x"77",   x"A9",   x"F6",   x"28",   x"89",   x"57", 
  x"37",   x"E9",   x"48",   x"96",   x"C9",   x"17",   x"B6",   x"68", 
  x"8A",   x"54",   x"F5",   x"2B",   x"74",   x"AA",   x"0B",   x"D5", 
  x"B5",   x"6B",   x"CA",   x"14",   x"4B",   x"95",   x"34",   x"EA", 
  x"F4",   x"2A",   x"8B",   x"55",   x"0A",   x"D4",   x"75",   x"AB", 
  x"CB",   x"15",   x"B4",   x"6A",   x"35",   x"EB",   x"4A",   x"94", 
  x"4D",   x"93",   x"32",   x"EC",   x"B3",   x"6D",   x"CC",   x"12", 
  x"72",   x"AC",   x"0D",   x"D3",   x"8C",   x"52",   x"F3",   x"2D", 
  x"33",   x"ED",   x"4C",   x"92",   x"CD",   x"13",   x"B2",   x"6C", 
  x"0C",   x"D2",   x"73",   x"AD",   x"F2",   x"2C",   x"8D",   x"53", 
  x"B1",   x"6F",   x"CE",   x"10",   x"4F",   x"91",   x"30",   x"EE", 
  x"8E",   x"50",   x"F1",   x"2F",   x"70",   x"AE",   x"0F",   x"D1", 
  x"CF",   x"11",   x"B0",   x"6E",   x"31",   x"EF",   x"4E",   x"90", 
  x"F0",   x"2E",   x"8F",   x"51",   x"0E",   x"D0",   x"71",   x"AF", 
  x"00",   x"DF",   x"7D",   x"A2",   x"FA",   x"25",   x"87",   x"58", 
  x"37",   x"E8",   x"4A",   x"95",   x"CD",   x"12",   x"B0",   x"6F", 
  x"6E",   x"B1",   x"13",   x"CC",   x"94",   x"4B",   x"E9",   x"36", 
  x"59",   x"86",   x"24",   x"FB",   x"A3",   x"7C",   x"DE",   x"01", 
  x"DC",   x"03",   x"A1",   x"7E",   x"26",   x"F9",   x"5B",   x"84", 
  x"EB",   x"34",   x"96",   x"49",   x"11",   x"CE",   x"6C",   x"B3", 
  x"B2",   x"6D",   x"CF",   x"10",   x"48",   x"97",   x"35",   x"EA", 
  x"85",   x"5A",   x"F8",   x"27",   x"7F",   x"A0",   x"02",   x"DD", 
  x"7B",   x"A4",   x"06",   x"D9",   x"81",   x"5E",   x"FC",   x"23", 
  x"4C",   x"93",   x"31",   x"EE",   x"B6",   x"69",   x"CB",   x"14", 
  x"15",   x"CA",   x"68",   x"B7",   x"EF",   x"30",   x"92",   x"4D", 
  x"22",   x"FD",   x"5F",   x"80",   x"D8",   x"07",   x"A5",   x"7A", 
  x"A7",   x"78",   x"DA",   x"05",   x"5D",   x"82",   x"20",   x"FF", 
  x"90",   x"4F",   x"ED",   x"32",   x"6A",   x"B5",   x"17",   x"C8", 
  x"C9",   x"16",   x"B4",   x"6B",   x"33",   x"EC",   x"4E",   x"91", 
  x"FE",   x"21",   x"83",   x"5C",   x"04",   x"DB",   x"79",   x"A6", 
  x"F6",   x"29",   x"8B",   x"54",   x"0C",   x"D3",   x"71",   x"AE", 
  x"C1",   x"1E",   x"BC",   x"63",   x"3B",   x"E4",   x"46",   x"99", 
  x"98",   x"47",   x"E5",   x"3A",   x"62",   x"BD",   x"1F",   x"C0", 
  x"AF",   x"70",   x"D2",   x"0D",   x"55",   x"8A",   x"28",   x"F7", 
  x"2A",   x"F5",   x"57",   x"88",   x"D0",   x"0F",   x"AD",   x"72", 
  x"1D",   x"C2",   x"60",   x"BF",   x"E7",   x"38",   x"9A",   x"45", 
  x"44",   x"9B",   x"39",   x"E6",   x"BE",   x"61",   x"C3",   x"1C", 
  x"73",   x"AC",   x"0E",   x"D1",   x"89",   x"56",   x"F4",   x"2B", 
  x"8D",   x"52",   x"F0",   x"2F",   x"77",   x"A8",   x"0A",   x"D5", 
  x"BA",   x"65",   x"C7",   x"18",   x"40",   x"9F",   x"3D",   x"E2", 
  x"E3",   x"3C",   x"9E",   x"41",   x"19",   x"C6",   x"64",   x"BB", 
  x"D4",   x"0B",   x"A9",   x"76",   x"2E",   x"F1",   x"53",   x"8C", 
  x"51",   x"8E",   x"2C",   x"F3",   x"AB",   x"74",   x"D6",   x"09", 
  x"66",   x"B9",   x"1B",   x"C4",   x"9C",   x"43",   x"E1",   x"3E", 
  x"3F",   x"E0",   x"42",   x"9D",   x"C5",   x"1A",   x"B8",   x"67", 
  x"08",   x"D7",   x"75",   x"AA",   x"F2",   x"2D",   x"8F",   x"50", 
  x"00",   x"E0",   x"03",   x"E3",   x"06",   x"E6",   x"05",   x"E5", 
  x"0C",   x"EC",   x"0F",   x"EF",   x"0A",   x"EA",   x"09",   x"E9", 
  x"18",   x"F8",   x"1B",   x"FB",   x"1E",   x"FE",   x"1D",   x"FD", 
  x"14",   x"F4",   x"17",   x"F7",   x"12",   x"F2",   x"11",   x"F1", 
  x"30",   x"D0",   x"33",   x"D3",   x"36",   x"D6",   x"35",   x"D5", 
  x"3C",   x"DC",   x"3F",   x"DF",   x"3A",   x"DA",   x"39",   x"D9", 
  x"28",   x"C8",   x"2B",   x"CB",   x"2E",   x"CE",   x"2D",   x"CD", 
  x"24",   x"C4",   x"27",   x"C7",   x"22",   x"C2",   x"21",   x"C1", 
  x"60",   x"80",   x"63",   x"83",   x"66",   x"86",   x"65",   x"85", 
  x"6C",   x"8C",   x"6F",   x"8F",   x"6A",   x"8A",   x"69",   x"89", 
  x"78",   x"98",   x"7B",   x"9B",   x"7E",   x"9E",   x"7D",   x"9D", 
  x"74",   x"94",   x"77",   x"97",   x"72",   x"92",   x"71",   x"91", 
  x"50",   x"B0",   x"53",   x"B3",   x"56",   x"B6",   x"55",   x"B5", 
  x"5C",   x"BC",   x"5F",   x"BF",   x"5A",   x"BA",   x"59",   x"B9", 
  x"48",   x"A8",   x"4B",   x"AB",   x"4E",   x"AE",   x"4D",   x"AD", 
  x"44",   x"A4",   x"47",   x"A7",   x"42",   x"A2",   x"41",   x"A1", 
  x"C0",   x"20",   x"C3",   x"23",   x"C6",   x"26",   x"C5",   x"25", 
  x"CC",   x"2C",   x"CF",   x"2F",   x"CA",   x"2A",   x"C9",   x"29", 
  x"D8",   x"38",   x"DB",   x"3B",   x"DE",   x"3E",   x"DD",   x"3D", 
  x"D4",   x"34",   x"D7",   x"37",   x"D2",   x"32",   x"D1",   x"31", 
  x"F0",   x"10",   x"F3",   x"13",   x"F6",   x"16",   x"F5",   x"15", 
  x"FC",   x"1C",   x"FF",   x"1F",   x"FA",   x"1A",   x"F9",   x"19", 
  x"E8",   x"08",   x"EB",   x"0B",   x"EE",   x"0E",   x"ED",   x"0D", 
  x"E4",   x"04",   x"E7",   x"07",   x"E2",   x"02",   x"E1",   x"01", 
  x"A0",   x"40",   x"A3",   x"43",   x"A6",   x"46",   x"A5",   x"45", 
  x"AC",   x"4C",   x"AF",   x"4F",   x"AA",   x"4A",   x"A9",   x"49", 
  x"B8",   x"58",   x"BB",   x"5B",   x"BE",   x"5E",   x"BD",   x"5D", 
  x"B4",   x"54",   x"B7",   x"57",   x"B2",   x"52",   x"B1",   x"51", 
  x"90",   x"70",   x"93",   x"73",   x"96",   x"76",   x"95",   x"75", 
  x"9C",   x"7C",   x"9F",   x"7F",   x"9A",   x"7A",   x"99",   x"79", 
  x"88",   x"68",   x"8B",   x"6B",   x"8E",   x"6E",   x"8D",   x"6D", 
  x"84",   x"64",   x"87",   x"67",   x"82",   x"62",   x"81",   x"61", 
  x"00",   x"E1",   x"01",   x"E0",   x"02",   x"E3",   x"03",   x"E2", 
  x"04",   x"E5",   x"05",   x"E4",   x"06",   x"E7",   x"07",   x"E6", 
  x"08",   x"E9",   x"09",   x"E8",   x"0A",   x"EB",   x"0B",   x"EA", 
  x"0C",   x"ED",   x"0D",   x"EC",   x"0E",   x"EF",   x"0F",   x"EE", 
  x"10",   x"F1",   x"11",   x"F0",   x"12",   x"F3",   x"13",   x"F2", 
  x"14",   x"F5",   x"15",   x"F4",   x"16",   x"F7",   x"17",   x"F6", 
  x"18",   x"F9",   x"19",   x"F8",   x"1A",   x"FB",   x"1B",   x"FA", 
  x"1C",   x"FD",   x"1D",   x"FC",   x"1E",   x"FF",   x"1F",   x"FE", 
  x"20",   x"C1",   x"21",   x"C0",   x"22",   x"C3",   x"23",   x"C2", 
  x"24",   x"C5",   x"25",   x"C4",   x"26",   x"C7",   x"27",   x"C6", 
  x"28",   x"C9",   x"29",   x"C8",   x"2A",   x"CB",   x"2B",   x"CA", 
  x"2C",   x"CD",   x"2D",   x"CC",   x"2E",   x"CF",   x"2F",   x"CE", 
  x"30",   x"D1",   x"31",   x"D0",   x"32",   x"D3",   x"33",   x"D2", 
  x"34",   x"D5",   x"35",   x"D4",   x"36",   x"D7",   x"37",   x"D6", 
  x"38",   x"D9",   x"39",   x"D8",   x"3A",   x"DB",   x"3B",   x"DA", 
  x"3C",   x"DD",   x"3D",   x"DC",   x"3E",   x"DF",   x"3F",   x"DE", 
  x"40",   x"A1",   x"41",   x"A0",   x"42",   x"A3",   x"43",   x"A2", 
  x"44",   x"A5",   x"45",   x"A4",   x"46",   x"A7",   x"47",   x"A6", 
  x"48",   x"A9",   x"49",   x"A8",   x"4A",   x"AB",   x"4B",   x"AA", 
  x"4C",   x"AD",   x"4D",   x"AC",   x"4E",   x"AF",   x"4F",   x"AE", 
  x"50",   x"B1",   x"51",   x"B0",   x"52",   x"B3",   x"53",   x"B2", 
  x"54",   x"B5",   x"55",   x"B4",   x"56",   x"B7",   x"57",   x"B6", 
  x"58",   x"B9",   x"59",   x"B8",   x"5A",   x"BB",   x"5B",   x"BA", 
  x"5C",   x"BD",   x"5D",   x"BC",   x"5E",   x"BF",   x"5F",   x"BE", 
  x"60",   x"81",   x"61",   x"80",   x"62",   x"83",   x"63",   x"82", 
  x"64",   x"85",   x"65",   x"84",   x"66",   x"87",   x"67",   x"86", 
  x"68",   x"89",   x"69",   x"88",   x"6A",   x"8B",   x"6B",   x"8A", 
  x"6C",   x"8D",   x"6D",   x"8C",   x"6E",   x"8F",   x"6F",   x"8E", 
  x"70",   x"91",   x"71",   x"90",   x"72",   x"93",   x"73",   x"92", 
  x"74",   x"95",   x"75",   x"94",   x"76",   x"97",   x"77",   x"96", 
  x"78",   x"99",   x"79",   x"98",   x"7A",   x"9B",   x"7B",   x"9A", 
  x"7C",   x"9D",   x"7D",   x"9C",   x"7E",   x"9F",   x"7F",   x"9E", 
  x"00",   x"E2",   x"07",   x"E5",   x"0E",   x"EC",   x"09",   x"EB", 
  x"1C",   x"FE",   x"1B",   x"F9",   x"12",   x"F0",   x"15",   x"F7", 
  x"38",   x"DA",   x"3F",   x"DD",   x"36",   x"D4",   x"31",   x"D3", 
  x"24",   x"C6",   x"23",   x"C1",   x"2A",   x"C8",   x"2D",   x"CF", 
  x"70",   x"92",   x"77",   x"95",   x"7E",   x"9C",   x"79",   x"9B", 
  x"6C",   x"8E",   x"6B",   x"89",   x"62",   x"80",   x"65",   x"87", 
  x"48",   x"AA",   x"4F",   x"AD",   x"46",   x"A4",   x"41",   x"A3", 
  x"54",   x"B6",   x"53",   x"B1",   x"5A",   x"B8",   x"5D",   x"BF", 
  x"E0",   x"02",   x"E7",   x"05",   x"EE",   x"0C",   x"E9",   x"0B", 
  x"FC",   x"1E",   x"FB",   x"19",   x"F2",   x"10",   x"F5",   x"17", 
  x"D8",   x"3A",   x"DF",   x"3D",   x"D6",   x"34",   x"D1",   x"33", 
  x"C4",   x"26",   x"C3",   x"21",   x"CA",   x"28",   x"CD",   x"2F", 
  x"90",   x"72",   x"97",   x"75",   x"9E",   x"7C",   x"99",   x"7B", 
  x"8C",   x"6E",   x"8B",   x"69",   x"82",   x"60",   x"85",   x"67", 
  x"A8",   x"4A",   x"AF",   x"4D",   x"A6",   x"44",   x"A1",   x"43", 
  x"B4",   x"56",   x"B3",   x"51",   x"BA",   x"58",   x"BD",   x"5F", 
  x"03",   x"E1",   x"04",   x"E6",   x"0D",   x"EF",   x"0A",   x"E8", 
  x"1F",   x"FD",   x"18",   x"FA",   x"11",   x"F3",   x"16",   x"F4", 
  x"3B",   x"D9",   x"3C",   x"DE",   x"35",   x"D7",   x"32",   x"D0", 
  x"27",   x"C5",   x"20",   x"C2",   x"29",   x"CB",   x"2E",   x"CC", 
  x"73",   x"91",   x"74",   x"96",   x"7D",   x"9F",   x"7A",   x"98", 
  x"6F",   x"8D",   x"68",   x"8A",   x"61",   x"83",   x"66",   x"84", 
  x"4B",   x"A9",   x"4C",   x"AE",   x"45",   x"A7",   x"42",   x"A0", 
  x"57",   x"B5",   x"50",   x"B2",   x"59",   x"BB",   x"5E",   x"BC", 
  x"E3",   x"01",   x"E4",   x"06",   x"ED",   x"0F",   x"EA",   x"08", 
  x"FF",   x"1D",   x"F8",   x"1A",   x"F1",   x"13",   x"F6",   x"14", 
  x"DB",   x"39",   x"DC",   x"3E",   x"D5",   x"37",   x"D2",   x"30", 
  x"C7",   x"25",   x"C0",   x"22",   x"C9",   x"2B",   x"CE",   x"2C", 
  x"93",   x"71",   x"94",   x"76",   x"9D",   x"7F",   x"9A",   x"78", 
  x"8F",   x"6D",   x"88",   x"6A",   x"81",   x"63",   x"86",   x"64", 
  x"AB",   x"49",   x"AC",   x"4E",   x"A5",   x"47",   x"A2",   x"40", 
  x"B7",   x"55",   x"B0",   x"52",   x"B9",   x"5B",   x"BE",   x"5C", 
  x"00",   x"E3",   x"05",   x"E6",   x"0A",   x"E9",   x"0F",   x"EC", 
  x"14",   x"F7",   x"11",   x"F2",   x"1E",   x"FD",   x"1B",   x"F8", 
  x"28",   x"CB",   x"2D",   x"CE",   x"22",   x"C1",   x"27",   x"C4", 
  x"3C",   x"DF",   x"39",   x"DA",   x"36",   x"D5",   x"33",   x"D0", 
  x"50",   x"B3",   x"55",   x"B6",   x"5A",   x"B9",   x"5F",   x"BC", 
  x"44",   x"A7",   x"41",   x"A2",   x"4E",   x"AD",   x"4B",   x"A8", 
  x"78",   x"9B",   x"7D",   x"9E",   x"72",   x"91",   x"77",   x"94", 
  x"6C",   x"8F",   x"69",   x"8A",   x"66",   x"85",   x"63",   x"80", 
  x"A0",   x"43",   x"A5",   x"46",   x"AA",   x"49",   x"AF",   x"4C", 
  x"B4",   x"57",   x"B1",   x"52",   x"BE",   x"5D",   x"BB",   x"58", 
  x"88",   x"6B",   x"8D",   x"6E",   x"82",   x"61",   x"87",   x"64", 
  x"9C",   x"7F",   x"99",   x"7A",   x"96",   x"75",   x"93",   x"70", 
  x"F0",   x"13",   x"F5",   x"16",   x"FA",   x"19",   x"FF",   x"1C", 
  x"E4",   x"07",   x"E1",   x"02",   x"EE",   x"0D",   x"EB",   x"08", 
  x"D8",   x"3B",   x"DD",   x"3E",   x"D2",   x"31",   x"D7",   x"34", 
  x"CC",   x"2F",   x"C9",   x"2A",   x"C6",   x"25",   x"C3",   x"20", 
  x"83",   x"60",   x"86",   x"65",   x"89",   x"6A",   x"8C",   x"6F", 
  x"97",   x"74",   x"92",   x"71",   x"9D",   x"7E",   x"98",   x"7B", 
  x"AB",   x"48",   x"AE",   x"4D",   x"A1",   x"42",   x"A4",   x"47", 
  x"BF",   x"5C",   x"BA",   x"59",   x"B5",   x"56",   x"B0",   x"53", 
  x"D3",   x"30",   x"D6",   x"35",   x"D9",   x"3A",   x"DC",   x"3F", 
  x"C7",   x"24",   x"C2",   x"21",   x"CD",   x"2E",   x"C8",   x"2B", 
  x"FB",   x"18",   x"FE",   x"1D",   x"F1",   x"12",   x"F4",   x"17", 
  x"EF",   x"0C",   x"EA",   x"09",   x"E5",   x"06",   x"E0",   x"03", 
  x"23",   x"C0",   x"26",   x"C5",   x"29",   x"CA",   x"2C",   x"CF", 
  x"37",   x"D4",   x"32",   x"D1",   x"3D",   x"DE",   x"38",   x"DB", 
  x"0B",   x"E8",   x"0E",   x"ED",   x"01",   x"E2",   x"04",   x"E7", 
  x"1F",   x"FC",   x"1A",   x"F9",   x"15",   x"F6",   x"10",   x"F3", 
  x"73",   x"90",   x"76",   x"95",   x"79",   x"9A",   x"7C",   x"9F", 
  x"67",   x"84",   x"62",   x"81",   x"6D",   x"8E",   x"68",   x"8B", 
  x"5B",   x"B8",   x"5E",   x"BD",   x"51",   x"B2",   x"54",   x"B7", 
  x"4F",   x"AC",   x"4A",   x"A9",   x"45",   x"A6",   x"40",   x"A3", 
  x"00",   x"E4",   x"0B",   x"EF",   x"16",   x"F2",   x"1D",   x"F9", 
  x"2C",   x"C8",   x"27",   x"C3",   x"3A",   x"DE",   x"31",   x"D5", 
  x"58",   x"BC",   x"53",   x"B7",   x"4E",   x"AA",   x"45",   x"A1", 
  x"74",   x"90",   x"7F",   x"9B",   x"62",   x"86",   x"69",   x"8D", 
  x"B0",   x"54",   x"BB",   x"5F",   x"A6",   x"42",   x"AD",   x"49", 
  x"9C",   x"78",   x"97",   x"73",   x"8A",   x"6E",   x"81",   x"65", 
  x"E8",   x"0C",   x"E3",   x"07",   x"FE",   x"1A",   x"F5",   x"11", 
  x"C4",   x"20",   x"CF",   x"2B",   x"D2",   x"36",   x"D9",   x"3D", 
  x"A3",   x"47",   x"A8",   x"4C",   x"B5",   x"51",   x"BE",   x"5A", 
  x"8F",   x"6B",   x"84",   x"60",   x"99",   x"7D",   x"92",   x"76", 
  x"FB",   x"1F",   x"F0",   x"14",   x"ED",   x"09",   x"E6",   x"02", 
  x"D7",   x"33",   x"DC",   x"38",   x"C1",   x"25",   x"CA",   x"2E", 
  x"13",   x"F7",   x"18",   x"FC",   x"05",   x"E1",   x"0E",   x"EA", 
  x"3F",   x"DB",   x"34",   x"D0",   x"29",   x"CD",   x"22",   x"C6", 
  x"4B",   x"AF",   x"40",   x"A4",   x"5D",   x"B9",   x"56",   x"B2", 
  x"67",   x"83",   x"6C",   x"88",   x"71",   x"95",   x"7A",   x"9E", 
  x"85",   x"61",   x"8E",   x"6A",   x"93",   x"77",   x"98",   x"7C", 
  x"A9",   x"4D",   x"A2",   x"46",   x"BF",   x"5B",   x"B4",   x"50", 
  x"DD",   x"39",   x"D6",   x"32",   x"CB",   x"2F",   x"C0",   x"24", 
  x"F1",   x"15",   x"FA",   x"1E",   x"E7",   x"03",   x"EC",   x"08", 
  x"35",   x"D1",   x"3E",   x"DA",   x"23",   x"C7",   x"28",   x"CC", 
  x"19",   x"FD",   x"12",   x"F6",   x"0F",   x"EB",   x"04",   x"E0", 
  x"6D",   x"89",   x"66",   x"82",   x"7B",   x"9F",   x"70",   x"94", 
  x"41",   x"A5",   x"4A",   x"AE",   x"57",   x"B3",   x"5C",   x"B8", 
  x"26",   x"C2",   x"2D",   x"C9",   x"30",   x"D4",   x"3B",   x"DF", 
  x"0A",   x"EE",   x"01",   x"E5",   x"1C",   x"F8",   x"17",   x"F3", 
  x"7E",   x"9A",   x"75",   x"91",   x"68",   x"8C",   x"63",   x"87", 
  x"52",   x"B6",   x"59",   x"BD",   x"44",   x"A0",   x"4F",   x"AB", 
  x"96",   x"72",   x"9D",   x"79",   x"80",   x"64",   x"8B",   x"6F", 
  x"BA",   x"5E",   x"B1",   x"55",   x"AC",   x"48",   x"A7",   x"43", 
  x"CE",   x"2A",   x"C5",   x"21",   x"D8",   x"3C",   x"D3",   x"37", 
  x"E2",   x"06",   x"E9",   x"0D",   x"F4",   x"10",   x"FF",   x"1B", 
  x"00",   x"E5",   x"09",   x"EC",   x"12",   x"F7",   x"1B",   x"FE", 
  x"24",   x"C1",   x"2D",   x"C8",   x"36",   x"D3",   x"3F",   x"DA", 
  x"48",   x"AD",   x"41",   x"A4",   x"5A",   x"BF",   x"53",   x"B6", 
  x"6C",   x"89",   x"65",   x"80",   x"7E",   x"9B",   x"77",   x"92", 
  x"90",   x"75",   x"99",   x"7C",   x"82",   x"67",   x"8B",   x"6E", 
  x"B4",   x"51",   x"BD",   x"58",   x"A6",   x"43",   x"AF",   x"4A", 
  x"D8",   x"3D",   x"D1",   x"34",   x"CA",   x"2F",   x"C3",   x"26", 
  x"FC",   x"19",   x"F5",   x"10",   x"EE",   x"0B",   x"E7",   x"02", 
  x"E3",   x"06",   x"EA",   x"0F",   x"F1",   x"14",   x"F8",   x"1D", 
  x"C7",   x"22",   x"CE",   x"2B",   x"D5",   x"30",   x"DC",   x"39", 
  x"AB",   x"4E",   x"A2",   x"47",   x"B9",   x"5C",   x"B0",   x"55", 
  x"8F",   x"6A",   x"86",   x"63",   x"9D",   x"78",   x"94",   x"71", 
  x"73",   x"96",   x"7A",   x"9F",   x"61",   x"84",   x"68",   x"8D", 
  x"57",   x"B2",   x"5E",   x"BB",   x"45",   x"A0",   x"4C",   x"A9", 
  x"3B",   x"DE",   x"32",   x"D7",   x"29",   x"CC",   x"20",   x"C5", 
  x"1F",   x"FA",   x"16",   x"F3",   x"0D",   x"E8",   x"04",   x"E1", 
  x"05",   x"E0",   x"0C",   x"E9",   x"17",   x"F2",   x"1E",   x"FB", 
  x"21",   x"C4",   x"28",   x"CD",   x"33",   x"D6",   x"3A",   x"DF", 
  x"4D",   x"A8",   x"44",   x"A1",   x"5F",   x"BA",   x"56",   x"B3", 
  x"69",   x"8C",   x"60",   x"85",   x"7B",   x"9E",   x"72",   x"97", 
  x"95",   x"70",   x"9C",   x"79",   x"87",   x"62",   x"8E",   x"6B", 
  x"B1",   x"54",   x"B8",   x"5D",   x"A3",   x"46",   x"AA",   x"4F", 
  x"DD",   x"38",   x"D4",   x"31",   x"CF",   x"2A",   x"C6",   x"23", 
  x"F9",   x"1C",   x"F0",   x"15",   x"EB",   x"0E",   x"E2",   x"07", 
  x"E6",   x"03",   x"EF",   x"0A",   x"F4",   x"11",   x"FD",   x"18", 
  x"C2",   x"27",   x"CB",   x"2E",   x"D0",   x"35",   x"D9",   x"3C", 
  x"AE",   x"4B",   x"A7",   x"42",   x"BC",   x"59",   x"B5",   x"50", 
  x"8A",   x"6F",   x"83",   x"66",   x"98",   x"7D",   x"91",   x"74", 
  x"76",   x"93",   x"7F",   x"9A",   x"64",   x"81",   x"6D",   x"88", 
  x"52",   x"B7",   x"5B",   x"BE",   x"40",   x"A5",   x"49",   x"AC", 
  x"3E",   x"DB",   x"37",   x"D2",   x"2C",   x"C9",   x"25",   x"C0", 
  x"1A",   x"FF",   x"13",   x"F6",   x"08",   x"ED",   x"01",   x"E4", 
  x"00",   x"E6",   x"0F",   x"E9",   x"1E",   x"F8",   x"11",   x"F7", 
  x"3C",   x"DA",   x"33",   x"D5",   x"22",   x"C4",   x"2D",   x"CB", 
  x"78",   x"9E",   x"77",   x"91",   x"66",   x"80",   x"69",   x"8F", 
  x"44",   x"A2",   x"4B",   x"AD",   x"5A",   x"BC",   x"55",   x"B3", 
  x"F0",   x"16",   x"FF",   x"19",   x"EE",   x"08",   x"E1",   x"07", 
  x"CC",   x"2A",   x"C3",   x"25",   x"D2",   x"34",   x"DD",   x"3B", 
  x"88",   x"6E",   x"87",   x"61",   x"96",   x"70",   x"99",   x"7F", 
  x"B4",   x"52",   x"BB",   x"5D",   x"AA",   x"4C",   x"A5",   x"43", 
  x"23",   x"C5",   x"2C",   x"CA",   x"3D",   x"DB",   x"32",   x"D4", 
  x"1F",   x"F9",   x"10",   x"F6",   x"01",   x"E7",   x"0E",   x"E8", 
  x"5B",   x"BD",   x"54",   x"B2",   x"45",   x"A3",   x"4A",   x"AC", 
  x"67",   x"81",   x"68",   x"8E",   x"79",   x"9F",   x"76",   x"90", 
  x"D3",   x"35",   x"DC",   x"3A",   x"CD",   x"2B",   x"C2",   x"24", 
  x"EF",   x"09",   x"E0",   x"06",   x"F1",   x"17",   x"FE",   x"18", 
  x"AB",   x"4D",   x"A4",   x"42",   x"B5",   x"53",   x"BA",   x"5C", 
  x"97",   x"71",   x"98",   x"7E",   x"89",   x"6F",   x"86",   x"60", 
  x"46",   x"A0",   x"49",   x"AF",   x"58",   x"BE",   x"57",   x"B1", 
  x"7A",   x"9C",   x"75",   x"93",   x"64",   x"82",   x"6B",   x"8D", 
  x"3E",   x"D8",   x"31",   x"D7",   x"20",   x"C6",   x"2F",   x"C9", 
  x"02",   x"E4",   x"0D",   x"EB",   x"1C",   x"FA",   x"13",   x"F5", 
  x"B6",   x"50",   x"B9",   x"5F",   x"A8",   x"4E",   x"A7",   x"41", 
  x"8A",   x"6C",   x"85",   x"63",   x"94",   x"72",   x"9B",   x"7D", 
  x"CE",   x"28",   x"C1",   x"27",   x"D0",   x"36",   x"DF",   x"39", 
  x"F2",   x"14",   x"FD",   x"1B",   x"EC",   x"0A",   x"E3",   x"05", 
  x"65",   x"83",   x"6A",   x"8C",   x"7B",   x"9D",   x"74",   x"92", 
  x"59",   x"BF",   x"56",   x"B0",   x"47",   x"A1",   x"48",   x"AE", 
  x"1D",   x"FB",   x"12",   x"F4",   x"03",   x"E5",   x"0C",   x"EA", 
  x"21",   x"C7",   x"2E",   x"C8",   x"3F",   x"D9",   x"30",   x"D6", 
  x"95",   x"73",   x"9A",   x"7C",   x"8B",   x"6D",   x"84",   x"62", 
  x"A9",   x"4F",   x"A6",   x"40",   x"B7",   x"51",   x"B8",   x"5E", 
  x"ED",   x"0B",   x"E2",   x"04",   x"F3",   x"15",   x"FC",   x"1A", 
  x"D1",   x"37",   x"DE",   x"38",   x"CF",   x"29",   x"C0",   x"26", 
  x"00",   x"E7",   x"0D",   x"EA",   x"1A",   x"FD",   x"17",   x"F0", 
  x"34",   x"D3",   x"39",   x"DE",   x"2E",   x"C9",   x"23",   x"C4", 
  x"68",   x"8F",   x"65",   x"82",   x"72",   x"95",   x"7F",   x"98", 
  x"5C",   x"BB",   x"51",   x"B6",   x"46",   x"A1",   x"4B",   x"AC", 
  x"D0",   x"37",   x"DD",   x"3A",   x"CA",   x"2D",   x"C7",   x"20", 
  x"E4",   x"03",   x"E9",   x"0E",   x"FE",   x"19",   x"F3",   x"14", 
  x"B8",   x"5F",   x"B5",   x"52",   x"A2",   x"45",   x"AF",   x"48", 
  x"8C",   x"6B",   x"81",   x"66",   x"96",   x"71",   x"9B",   x"7C", 
  x"63",   x"84",   x"6E",   x"89",   x"79",   x"9E",   x"74",   x"93", 
  x"57",   x"B0",   x"5A",   x"BD",   x"4D",   x"AA",   x"40",   x"A7", 
  x"0B",   x"EC",   x"06",   x"E1",   x"11",   x"F6",   x"1C",   x"FB", 
  x"3F",   x"D8",   x"32",   x"D5",   x"25",   x"C2",   x"28",   x"CF", 
  x"B3",   x"54",   x"BE",   x"59",   x"A9",   x"4E",   x"A4",   x"43", 
  x"87",   x"60",   x"8A",   x"6D",   x"9D",   x"7A",   x"90",   x"77", 
  x"DB",   x"3C",   x"D6",   x"31",   x"C1",   x"26",   x"CC",   x"2B", 
  x"EF",   x"08",   x"E2",   x"05",   x"F5",   x"12",   x"F8",   x"1F", 
  x"C6",   x"21",   x"CB",   x"2C",   x"DC",   x"3B",   x"D1",   x"36", 
  x"F2",   x"15",   x"FF",   x"18",   x"E8",   x"0F",   x"E5",   x"02", 
  x"AE",   x"49",   x"A3",   x"44",   x"B4",   x"53",   x"B9",   x"5E", 
  x"9A",   x"7D",   x"97",   x"70",   x"80",   x"67",   x"8D",   x"6A", 
  x"16",   x"F1",   x"1B",   x"FC",   x"0C",   x"EB",   x"01",   x"E6", 
  x"22",   x"C5",   x"2F",   x"C8",   x"38",   x"DF",   x"35",   x"D2", 
  x"7E",   x"99",   x"73",   x"94",   x"64",   x"83",   x"69",   x"8E", 
  x"4A",   x"AD",   x"47",   x"A0",   x"50",   x"B7",   x"5D",   x"BA", 
  x"A5",   x"42",   x"A8",   x"4F",   x"BF",   x"58",   x"B2",   x"55", 
  x"91",   x"76",   x"9C",   x"7B",   x"8B",   x"6C",   x"86",   x"61", 
  x"CD",   x"2A",   x"C0",   x"27",   x"D7",   x"30",   x"DA",   x"3D", 
  x"F9",   x"1E",   x"F4",   x"13",   x"E3",   x"04",   x"EE",   x"09", 
  x"75",   x"92",   x"78",   x"9F",   x"6F",   x"88",   x"62",   x"85", 
  x"41",   x"A6",   x"4C",   x"AB",   x"5B",   x"BC",   x"56",   x"B1", 
  x"1D",   x"FA",   x"10",   x"F7",   x"07",   x"E0",   x"0A",   x"ED", 
  x"29",   x"CE",   x"24",   x"C3",   x"33",   x"D4",   x"3E",   x"D9", 
  x"00",   x"E8",   x"13",   x"FB",   x"26",   x"CE",   x"35",   x"DD", 
  x"4C",   x"A4",   x"5F",   x"B7",   x"6A",   x"82",   x"79",   x"91", 
  x"98",   x"70",   x"8B",   x"63",   x"BE",   x"56",   x"AD",   x"45", 
  x"D4",   x"3C",   x"C7",   x"2F",   x"F2",   x"1A",   x"E1",   x"09", 
  x"F3",   x"1B",   x"E0",   x"08",   x"D5",   x"3D",   x"C6",   x"2E", 
  x"BF",   x"57",   x"AC",   x"44",   x"99",   x"71",   x"8A",   x"62", 
  x"6B",   x"83",   x"78",   x"90",   x"4D",   x"A5",   x"5E",   x"B6", 
  x"27",   x"CF",   x"34",   x"DC",   x"01",   x"E9",   x"12",   x"FA", 
  x"25",   x"CD",   x"36",   x"DE",   x"03",   x"EB",   x"10",   x"F8", 
  x"69",   x"81",   x"7A",   x"92",   x"4F",   x"A7",   x"5C",   x"B4", 
  x"BD",   x"55",   x"AE",   x"46",   x"9B",   x"73",   x"88",   x"60", 
  x"F1",   x"19",   x"E2",   x"0A",   x"D7",   x"3F",   x"C4",   x"2C", 
  x"D6",   x"3E",   x"C5",   x"2D",   x"F0",   x"18",   x"E3",   x"0B", 
  x"9A",   x"72",   x"89",   x"61",   x"BC",   x"54",   x"AF",   x"47", 
  x"4E",   x"A6",   x"5D",   x"B5",   x"68",   x"80",   x"7B",   x"93", 
  x"02",   x"EA",   x"11",   x"F9",   x"24",   x"CC",   x"37",   x"DF", 
  x"4A",   x"A2",   x"59",   x"B1",   x"6C",   x"84",   x"7F",   x"97", 
  x"06",   x"EE",   x"15",   x"FD",   x"20",   x"C8",   x"33",   x"DB", 
  x"D2",   x"3A",   x"C1",   x"29",   x"F4",   x"1C",   x"E7",   x"0F", 
  x"9E",   x"76",   x"8D",   x"65",   x"B8",   x"50",   x"AB",   x"43", 
  x"B9",   x"51",   x"AA",   x"42",   x"9F",   x"77",   x"8C",   x"64", 
  x"F5",   x"1D",   x"E6",   x"0E",   x"D3",   x"3B",   x"C0",   x"28", 
  x"21",   x"C9",   x"32",   x"DA",   x"07",   x"EF",   x"14",   x"FC", 
  x"6D",   x"85",   x"7E",   x"96",   x"4B",   x"A3",   x"58",   x"B0", 
  x"6F",   x"87",   x"7C",   x"94",   x"49",   x"A1",   x"5A",   x"B2", 
  x"23",   x"CB",   x"30",   x"D8",   x"05",   x"ED",   x"16",   x"FE", 
  x"F7",   x"1F",   x"E4",   x"0C",   x"D1",   x"39",   x"C2",   x"2A", 
  x"BB",   x"53",   x"A8",   x"40",   x"9D",   x"75",   x"8E",   x"66", 
  x"9C",   x"74",   x"8F",   x"67",   x"BA",   x"52",   x"A9",   x"41", 
  x"D0",   x"38",   x"C3",   x"2B",   x"F6",   x"1E",   x"E5",   x"0D", 
  x"04",   x"EC",   x"17",   x"FF",   x"22",   x"CA",   x"31",   x"D9", 
  x"48",   x"A0",   x"5B",   x"B3",   x"6E",   x"86",   x"7D",   x"95", 
  x"00",   x"E9",   x"11",   x"F8",   x"22",   x"CB",   x"33",   x"DA", 
  x"44",   x"AD",   x"55",   x"BC",   x"66",   x"8F",   x"77",   x"9E", 
  x"88",   x"61",   x"99",   x"70",   x"AA",   x"43",   x"BB",   x"52", 
  x"CC",   x"25",   x"DD",   x"34",   x"EE",   x"07",   x"FF",   x"16", 
  x"D3",   x"3A",   x"C2",   x"2B",   x"F1",   x"18",   x"E0",   x"09", 
  x"97",   x"7E",   x"86",   x"6F",   x"B5",   x"5C",   x"A4",   x"4D", 
  x"5B",   x"B2",   x"4A",   x"A3",   x"79",   x"90",   x"68",   x"81", 
  x"1F",   x"F6",   x"0E",   x"E7",   x"3D",   x"D4",   x"2C",   x"C5", 
  x"65",   x"8C",   x"74",   x"9D",   x"47",   x"AE",   x"56",   x"BF", 
  x"21",   x"C8",   x"30",   x"D9",   x"03",   x"EA",   x"12",   x"FB", 
  x"ED",   x"04",   x"FC",   x"15",   x"CF",   x"26",   x"DE",   x"37", 
  x"A9",   x"40",   x"B8",   x"51",   x"8B",   x"62",   x"9A",   x"73", 
  x"B6",   x"5F",   x"A7",   x"4E",   x"94",   x"7D",   x"85",   x"6C", 
  x"F2",   x"1B",   x"E3",   x"0A",   x"D0",   x"39",   x"C1",   x"28", 
  x"3E",   x"D7",   x"2F",   x"C6",   x"1C",   x"F5",   x"0D",   x"E4", 
  x"7A",   x"93",   x"6B",   x"82",   x"58",   x"B1",   x"49",   x"A0", 
  x"CA",   x"23",   x"DB",   x"32",   x"E8",   x"01",   x"F9",   x"10", 
  x"8E",   x"67",   x"9F",   x"76",   x"AC",   x"45",   x"BD",   x"54", 
  x"42",   x"AB",   x"53",   x"BA",   x"60",   x"89",   x"71",   x"98", 
  x"06",   x"EF",   x"17",   x"FE",   x"24",   x"CD",   x"35",   x"DC", 
  x"19",   x"F0",   x"08",   x"E1",   x"3B",   x"D2",   x"2A",   x"C3", 
  x"5D",   x"B4",   x"4C",   x"A5",   x"7F",   x"96",   x"6E",   x"87", 
  x"91",   x"78",   x"80",   x"69",   x"B3",   x"5A",   x"A2",   x"4B", 
  x"D5",   x"3C",   x"C4",   x"2D",   x"F7",   x"1E",   x"E6",   x"0F", 
  x"AF",   x"46",   x"BE",   x"57",   x"8D",   x"64",   x"9C",   x"75", 
  x"EB",   x"02",   x"FA",   x"13",   x"C9",   x"20",   x"D8",   x"31", 
  x"27",   x"CE",   x"36",   x"DF",   x"05",   x"EC",   x"14",   x"FD", 
  x"63",   x"8A",   x"72",   x"9B",   x"41",   x"A8",   x"50",   x"B9", 
  x"7C",   x"95",   x"6D",   x"84",   x"5E",   x"B7",   x"4F",   x"A6", 
  x"38",   x"D1",   x"29",   x"C0",   x"1A",   x"F3",   x"0B",   x"E2", 
  x"F4",   x"1D",   x"E5",   x"0C",   x"D6",   x"3F",   x"C7",   x"2E", 
  x"B0",   x"59",   x"A1",   x"48",   x"92",   x"7B",   x"83",   x"6A", 
  x"00",   x"EA",   x"17",   x"FD",   x"2E",   x"C4",   x"39",   x"D3", 
  x"5C",   x"B6",   x"4B",   x"A1",   x"72",   x"98",   x"65",   x"8F", 
  x"B8",   x"52",   x"AF",   x"45",   x"96",   x"7C",   x"81",   x"6B", 
  x"E4",   x"0E",   x"F3",   x"19",   x"CA",   x"20",   x"DD",   x"37", 
  x"B3",   x"59",   x"A4",   x"4E",   x"9D",   x"77",   x"8A",   x"60", 
  x"EF",   x"05",   x"F8",   x"12",   x"C1",   x"2B",   x"D6",   x"3C", 
  x"0B",   x"E1",   x"1C",   x"F6",   x"25",   x"CF",   x"32",   x"D8", 
  x"57",   x"BD",   x"40",   x"AA",   x"79",   x"93",   x"6E",   x"84", 
  x"A5",   x"4F",   x"B2",   x"58",   x"8B",   x"61",   x"9C",   x"76", 
  x"F9",   x"13",   x"EE",   x"04",   x"D7",   x"3D",   x"C0",   x"2A", 
  x"1D",   x"F7",   x"0A",   x"E0",   x"33",   x"D9",   x"24",   x"CE", 
  x"41",   x"AB",   x"56",   x"BC",   x"6F",   x"85",   x"78",   x"92", 
  x"16",   x"FC",   x"01",   x"EB",   x"38",   x"D2",   x"2F",   x"C5", 
  x"4A",   x"A0",   x"5D",   x"B7",   x"64",   x"8E",   x"73",   x"99", 
  x"AE",   x"44",   x"B9",   x"53",   x"80",   x"6A",   x"97",   x"7D", 
  x"F2",   x"18",   x"E5",   x"0F",   x"DC",   x"36",   x"CB",   x"21", 
  x"89",   x"63",   x"9E",   x"74",   x"A7",   x"4D",   x"B0",   x"5A", 
  x"D5",   x"3F",   x"C2",   x"28",   x"FB",   x"11",   x"EC",   x"06", 
  x"31",   x"DB",   x"26",   x"CC",   x"1F",   x"F5",   x"08",   x"E2", 
  x"6D",   x"87",   x"7A",   x"90",   x"43",   x"A9",   x"54",   x"BE", 
  x"3A",   x"D0",   x"2D",   x"C7",   x"14",   x"FE",   x"03",   x"E9", 
  x"66",   x"8C",   x"71",   x"9B",   x"48",   x"A2",   x"5F",   x"B5", 
  x"82",   x"68",   x"95",   x"7F",   x"AC",   x"46",   x"BB",   x"51", 
  x"DE",   x"34",   x"C9",   x"23",   x"F0",   x"1A",   x"E7",   x"0D", 
  x"2C",   x"C6",   x"3B",   x"D1",   x"02",   x"E8",   x"15",   x"FF", 
  x"70",   x"9A",   x"67",   x"8D",   x"5E",   x"B4",   x"49",   x"A3", 
  x"94",   x"7E",   x"83",   x"69",   x"BA",   x"50",   x"AD",   x"47", 
  x"C8",   x"22",   x"DF",   x"35",   x"E6",   x"0C",   x"F1",   x"1B", 
  x"9F",   x"75",   x"88",   x"62",   x"B1",   x"5B",   x"A6",   x"4C", 
  x"C3",   x"29",   x"D4",   x"3E",   x"ED",   x"07",   x"FA",   x"10", 
  x"27",   x"CD",   x"30",   x"DA",   x"09",   x"E3",   x"1E",   x"F4", 
  x"7B",   x"91",   x"6C",   x"86",   x"55",   x"BF",   x"42",   x"A8", 
  x"00",   x"EB",   x"15",   x"FE",   x"2A",   x"C1",   x"3F",   x"D4", 
  x"54",   x"BF",   x"41",   x"AA",   x"7E",   x"95",   x"6B",   x"80", 
  x"A8",   x"43",   x"BD",   x"56",   x"82",   x"69",   x"97",   x"7C", 
  x"FC",   x"17",   x"E9",   x"02",   x"D6",   x"3D",   x"C3",   x"28", 
  x"93",   x"78",   x"86",   x"6D",   x"B9",   x"52",   x"AC",   x"47", 
  x"C7",   x"2C",   x"D2",   x"39",   x"ED",   x"06",   x"F8",   x"13", 
  x"3B",   x"D0",   x"2E",   x"C5",   x"11",   x"FA",   x"04",   x"EF", 
  x"6F",   x"84",   x"7A",   x"91",   x"45",   x"AE",   x"50",   x"BB", 
  x"E5",   x"0E",   x"F0",   x"1B",   x"CF",   x"24",   x"DA",   x"31", 
  x"B1",   x"5A",   x"A4",   x"4F",   x"9B",   x"70",   x"8E",   x"65", 
  x"4D",   x"A6",   x"58",   x"B3",   x"67",   x"8C",   x"72",   x"99", 
  x"19",   x"F2",   x"0C",   x"E7",   x"33",   x"D8",   x"26",   x"CD", 
  x"76",   x"9D",   x"63",   x"88",   x"5C",   x"B7",   x"49",   x"A2", 
  x"22",   x"C9",   x"37",   x"DC",   x"08",   x"E3",   x"1D",   x"F6", 
  x"DE",   x"35",   x"CB",   x"20",   x"F4",   x"1F",   x"E1",   x"0A", 
  x"8A",   x"61",   x"9F",   x"74",   x"A0",   x"4B",   x"B5",   x"5E", 
  x"09",   x"E2",   x"1C",   x"F7",   x"23",   x"C8",   x"36",   x"DD", 
  x"5D",   x"B6",   x"48",   x"A3",   x"77",   x"9C",   x"62",   x"89", 
  x"A1",   x"4A",   x"B4",   x"5F",   x"8B",   x"60",   x"9E",   x"75", 
  x"F5",   x"1E",   x"E0",   x"0B",   x"DF",   x"34",   x"CA",   x"21", 
  x"9A",   x"71",   x"8F",   x"64",   x"B0",   x"5B",   x"A5",   x"4E", 
  x"CE",   x"25",   x"DB",   x"30",   x"E4",   x"0F",   x"F1",   x"1A", 
  x"32",   x"D9",   x"27",   x"CC",   x"18",   x"F3",   x"0D",   x"E6", 
  x"66",   x"8D",   x"73",   x"98",   x"4C",   x"A7",   x"59",   x"B2", 
  x"EC",   x"07",   x"F9",   x"12",   x"C6",   x"2D",   x"D3",   x"38", 
  x"B8",   x"53",   x"AD",   x"46",   x"92",   x"79",   x"87",   x"6C", 
  x"44",   x"AF",   x"51",   x"BA",   x"6E",   x"85",   x"7B",   x"90", 
  x"10",   x"FB",   x"05",   x"EE",   x"3A",   x"D1",   x"2F",   x"C4", 
  x"7F",   x"94",   x"6A",   x"81",   x"55",   x"BE",   x"40",   x"AB", 
  x"2B",   x"C0",   x"3E",   x"D5",   x"01",   x"EA",   x"14",   x"FF", 
  x"D7",   x"3C",   x"C2",   x"29",   x"FD",   x"16",   x"E8",   x"03", 
  x"83",   x"68",   x"96",   x"7D",   x"A9",   x"42",   x"BC",   x"57", 
  x"00",   x"EC",   x"1B",   x"F7",   x"36",   x"DA",   x"2D",   x"C1", 
  x"6C",   x"80",   x"77",   x"9B",   x"5A",   x"B6",   x"41",   x"AD", 
  x"D8",   x"34",   x"C3",   x"2F",   x"EE",   x"02",   x"F5",   x"19", 
  x"B4",   x"58",   x"AF",   x"43",   x"82",   x"6E",   x"99",   x"75", 
  x"73",   x"9F",   x"68",   x"84",   x"45",   x"A9",   x"5E",   x"B2", 
  x"1F",   x"F3",   x"04",   x"E8",   x"29",   x"C5",   x"32",   x"DE", 
  x"AB",   x"47",   x"B0",   x"5C",   x"9D",   x"71",   x"86",   x"6A", 
  x"C7",   x"2B",   x"DC",   x"30",   x"F1",   x"1D",   x"EA",   x"06", 
  x"E6",   x"0A",   x"FD",   x"11",   x"D0",   x"3C",   x"CB",   x"27", 
  x"8A",   x"66",   x"91",   x"7D",   x"BC",   x"50",   x"A7",   x"4B", 
  x"3E",   x"D2",   x"25",   x"C9",   x"08",   x"E4",   x"13",   x"FF", 
  x"52",   x"BE",   x"49",   x"A5",   x"64",   x"88",   x"7F",   x"93", 
  x"95",   x"79",   x"8E",   x"62",   x"A3",   x"4F",   x"B8",   x"54", 
  x"F9",   x"15",   x"E2",   x"0E",   x"CF",   x"23",   x"D4",   x"38", 
  x"4D",   x"A1",   x"56",   x"BA",   x"7B",   x"97",   x"60",   x"8C", 
  x"21",   x"CD",   x"3A",   x"D6",   x"17",   x"FB",   x"0C",   x"E0", 
  x"0F",   x"E3",   x"14",   x"F8",   x"39",   x"D5",   x"22",   x"CE", 
  x"63",   x"8F",   x"78",   x"94",   x"55",   x"B9",   x"4E",   x"A2", 
  x"D7",   x"3B",   x"CC",   x"20",   x"E1",   x"0D",   x"FA",   x"16", 
  x"BB",   x"57",   x"A0",   x"4C",   x"8D",   x"61",   x"96",   x"7A", 
  x"7C",   x"90",   x"67",   x"8B",   x"4A",   x"A6",   x"51",   x"BD", 
  x"10",   x"FC",   x"0B",   x"E7",   x"26",   x"CA",   x"3D",   x"D1", 
  x"A4",   x"48",   x"BF",   x"53",   x"92",   x"7E",   x"89",   x"65", 
  x"C8",   x"24",   x"D3",   x"3F",   x"FE",   x"12",   x"E5",   x"09", 
  x"E9",   x"05",   x"F2",   x"1E",   x"DF",   x"33",   x"C4",   x"28", 
  x"85",   x"69",   x"9E",   x"72",   x"B3",   x"5F",   x"A8",   x"44", 
  x"31",   x"DD",   x"2A",   x"C6",   x"07",   x"EB",   x"1C",   x"F0", 
  x"5D",   x"B1",   x"46",   x"AA",   x"6B",   x"87",   x"70",   x"9C", 
  x"9A",   x"76",   x"81",   x"6D",   x"AC",   x"40",   x"B7",   x"5B", 
  x"F6",   x"1A",   x"ED",   x"01",   x"C0",   x"2C",   x"DB",   x"37", 
  x"42",   x"AE",   x"59",   x"B5",   x"74",   x"98",   x"6F",   x"83", 
  x"2E",   x"C2",   x"35",   x"D9",   x"18",   x"F4",   x"03",   x"EF", 
  x"00",   x"ED",   x"19",   x"F4",   x"32",   x"DF",   x"2B",   x"C6", 
  x"64",   x"89",   x"7D",   x"90",   x"56",   x"BB",   x"4F",   x"A2", 
  x"C8",   x"25",   x"D1",   x"3C",   x"FA",   x"17",   x"E3",   x"0E", 
  x"AC",   x"41",   x"B5",   x"58",   x"9E",   x"73",   x"87",   x"6A", 
  x"53",   x"BE",   x"4A",   x"A7",   x"61",   x"8C",   x"78",   x"95", 
  x"37",   x"DA",   x"2E",   x"C3",   x"05",   x"E8",   x"1C",   x"F1", 
  x"9B",   x"76",   x"82",   x"6F",   x"A9",   x"44",   x"B0",   x"5D", 
  x"FF",   x"12",   x"E6",   x"0B",   x"CD",   x"20",   x"D4",   x"39", 
  x"A6",   x"4B",   x"BF",   x"52",   x"94",   x"79",   x"8D",   x"60", 
  x"C2",   x"2F",   x"DB",   x"36",   x"F0",   x"1D",   x"E9",   x"04", 
  x"6E",   x"83",   x"77",   x"9A",   x"5C",   x"B1",   x"45",   x"A8", 
  x"0A",   x"E7",   x"13",   x"FE",   x"38",   x"D5",   x"21",   x"CC", 
  x"F5",   x"18",   x"EC",   x"01",   x"C7",   x"2A",   x"DE",   x"33", 
  x"91",   x"7C",   x"88",   x"65",   x"A3",   x"4E",   x"BA",   x"57", 
  x"3D",   x"D0",   x"24",   x"C9",   x"0F",   x"E2",   x"16",   x"FB", 
  x"59",   x"B4",   x"40",   x"AD",   x"6B",   x"86",   x"72",   x"9F", 
  x"8F",   x"62",   x"96",   x"7B",   x"BD",   x"50",   x"A4",   x"49", 
  x"EB",   x"06",   x"F2",   x"1F",   x"D9",   x"34",   x"C0",   x"2D", 
  x"47",   x"AA",   x"5E",   x"B3",   x"75",   x"98",   x"6C",   x"81", 
  x"23",   x"CE",   x"3A",   x"D7",   x"11",   x"FC",   x"08",   x"E5", 
  x"DC",   x"31",   x"C5",   x"28",   x"EE",   x"03",   x"F7",   x"1A", 
  x"B8",   x"55",   x"A1",   x"4C",   x"8A",   x"67",   x"93",   x"7E", 
  x"14",   x"F9",   x"0D",   x"E0",   x"26",   x"CB",   x"3F",   x"D2", 
  x"70",   x"9D",   x"69",   x"84",   x"42",   x"AF",   x"5B",   x"B6", 
  x"29",   x"C4",   x"30",   x"DD",   x"1B",   x"F6",   x"02",   x"EF", 
  x"4D",   x"A0",   x"54",   x"B9",   x"7F",   x"92",   x"66",   x"8B", 
  x"E1",   x"0C",   x"F8",   x"15",   x"D3",   x"3E",   x"CA",   x"27", 
  x"85",   x"68",   x"9C",   x"71",   x"B7",   x"5A",   x"AE",   x"43", 
  x"7A",   x"97",   x"63",   x"8E",   x"48",   x"A5",   x"51",   x"BC", 
  x"1E",   x"F3",   x"07",   x"EA",   x"2C",   x"C1",   x"35",   x"D8", 
  x"B2",   x"5F",   x"AB",   x"46",   x"80",   x"6D",   x"99",   x"74", 
  x"D6",   x"3B",   x"CF",   x"22",   x"E4",   x"09",   x"FD",   x"10", 
  x"00",   x"EE",   x"1F",   x"F1",   x"3E",   x"D0",   x"21",   x"CF", 
  x"7C",   x"92",   x"63",   x"8D",   x"42",   x"AC",   x"5D",   x"B3", 
  x"F8",   x"16",   x"E7",   x"09",   x"C6",   x"28",   x"D9",   x"37", 
  x"84",   x"6A",   x"9B",   x"75",   x"BA",   x"54",   x"A5",   x"4B", 
  x"33",   x"DD",   x"2C",   x"C2",   x"0D",   x"E3",   x"12",   x"FC", 
  x"4F",   x"A1",   x"50",   x"BE",   x"71",   x"9F",   x"6E",   x"80", 
  x"CB",   x"25",   x"D4",   x"3A",   x"F5",   x"1B",   x"EA",   x"04", 
  x"B7",   x"59",   x"A8",   x"46",   x"89",   x"67",   x"96",   x"78", 
  x"66",   x"88",   x"79",   x"97",   x"58",   x"B6",   x"47",   x"A9", 
  x"1A",   x"F4",   x"05",   x"EB",   x"24",   x"CA",   x"3B",   x"D5", 
  x"9E",   x"70",   x"81",   x"6F",   x"A0",   x"4E",   x"BF",   x"51", 
  x"E2",   x"0C",   x"FD",   x"13",   x"DC",   x"32",   x"C3",   x"2D", 
  x"55",   x"BB",   x"4A",   x"A4",   x"6B",   x"85",   x"74",   x"9A", 
  x"29",   x"C7",   x"36",   x"D8",   x"17",   x"F9",   x"08",   x"E6", 
  x"AD",   x"43",   x"B2",   x"5C",   x"93",   x"7D",   x"8C",   x"62", 
  x"D1",   x"3F",   x"CE",   x"20",   x"EF",   x"01",   x"F0",   x"1E", 
  x"CC",   x"22",   x"D3",   x"3D",   x"F2",   x"1C",   x"ED",   x"03", 
  x"B0",   x"5E",   x"AF",   x"41",   x"8E",   x"60",   x"91",   x"7F", 
  x"34",   x"DA",   x"2B",   x"C5",   x"0A",   x"E4",   x"15",   x"FB", 
  x"48",   x"A6",   x"57",   x"B9",   x"76",   x"98",   x"69",   x"87", 
  x"FF",   x"11",   x"E0",   x"0E",   x"C1",   x"2F",   x"DE",   x"30", 
  x"83",   x"6D",   x"9C",   x"72",   x"BD",   x"53",   x"A2",   x"4C", 
  x"07",   x"E9",   x"18",   x"F6",   x"39",   x"D7",   x"26",   x"C8", 
  x"7B",   x"95",   x"64",   x"8A",   x"45",   x"AB",   x"5A",   x"B4", 
  x"AA",   x"44",   x"B5",   x"5B",   x"94",   x"7A",   x"8B",   x"65", 
  x"D6",   x"38",   x"C9",   x"27",   x"E8",   x"06",   x"F7",   x"19", 
  x"52",   x"BC",   x"4D",   x"A3",   x"6C",   x"82",   x"73",   x"9D", 
  x"2E",   x"C0",   x"31",   x"DF",   x"10",   x"FE",   x"0F",   x"E1", 
  x"99",   x"77",   x"86",   x"68",   x"A7",   x"49",   x"B8",   x"56", 
  x"E5",   x"0B",   x"FA",   x"14",   x"DB",   x"35",   x"C4",   x"2A", 
  x"61",   x"8F",   x"7E",   x"90",   x"5F",   x"B1",   x"40",   x"AE", 
  x"1D",   x"F3",   x"02",   x"EC",   x"23",   x"CD",   x"3C",   x"D2", 
  x"00",   x"EF",   x"1D",   x"F2",   x"3A",   x"D5",   x"27",   x"C8", 
  x"74",   x"9B",   x"69",   x"86",   x"4E",   x"A1",   x"53",   x"BC", 
  x"E8",   x"07",   x"F5",   x"1A",   x"D2",   x"3D",   x"CF",   x"20", 
  x"9C",   x"73",   x"81",   x"6E",   x"A6",   x"49",   x"BB",   x"54", 
  x"13",   x"FC",   x"0E",   x"E1",   x"29",   x"C6",   x"34",   x"DB", 
  x"67",   x"88",   x"7A",   x"95",   x"5D",   x"B2",   x"40",   x"AF", 
  x"FB",   x"14",   x"E6",   x"09",   x"C1",   x"2E",   x"DC",   x"33", 
  x"8F",   x"60",   x"92",   x"7D",   x"B5",   x"5A",   x"A8",   x"47", 
  x"26",   x"C9",   x"3B",   x"D4",   x"1C",   x"F3",   x"01",   x"EE", 
  x"52",   x"BD",   x"4F",   x"A0",   x"68",   x"87",   x"75",   x"9A", 
  x"CE",   x"21",   x"D3",   x"3C",   x"F4",   x"1B",   x"E9",   x"06", 
  x"BA",   x"55",   x"A7",   x"48",   x"80",   x"6F",   x"9D",   x"72", 
  x"35",   x"DA",   x"28",   x"C7",   x"0F",   x"E0",   x"12",   x"FD", 
  x"41",   x"AE",   x"5C",   x"B3",   x"7B",   x"94",   x"66",   x"89", 
  x"DD",   x"32",   x"C0",   x"2F",   x"E7",   x"08",   x"FA",   x"15", 
  x"A9",   x"46",   x"B4",   x"5B",   x"93",   x"7C",   x"8E",   x"61", 
  x"4C",   x"A3",   x"51",   x"BE",   x"76",   x"99",   x"6B",   x"84", 
  x"38",   x"D7",   x"25",   x"CA",   x"02",   x"ED",   x"1F",   x"F0", 
  x"A4",   x"4B",   x"B9",   x"56",   x"9E",   x"71",   x"83",   x"6C", 
  x"D0",   x"3F",   x"CD",   x"22",   x"EA",   x"05",   x"F7",   x"18", 
  x"5F",   x"B0",   x"42",   x"AD",   x"65",   x"8A",   x"78",   x"97", 
  x"2B",   x"C4",   x"36",   x"D9",   x"11",   x"FE",   x"0C",   x"E3", 
  x"B7",   x"58",   x"AA",   x"45",   x"8D",   x"62",   x"90",   x"7F", 
  x"C3",   x"2C",   x"DE",   x"31",   x"F9",   x"16",   x"E4",   x"0B", 
  x"6A",   x"85",   x"77",   x"98",   x"50",   x"BF",   x"4D",   x"A2", 
  x"1E",   x"F1",   x"03",   x"EC",   x"24",   x"CB",   x"39",   x"D6", 
  x"82",   x"6D",   x"9F",   x"70",   x"B8",   x"57",   x"A5",   x"4A", 
  x"F6",   x"19",   x"EB",   x"04",   x"CC",   x"23",   x"D1",   x"3E", 
  x"79",   x"96",   x"64",   x"8B",   x"43",   x"AC",   x"5E",   x"B1", 
  x"0D",   x"E2",   x"10",   x"FF",   x"37",   x"D8",   x"2A",   x"C5", 
  x"91",   x"7E",   x"8C",   x"63",   x"AB",   x"44",   x"B6",   x"59", 
  x"E5",   x"0A",   x"F8",   x"17",   x"DF",   x"30",   x"C2",   x"2D", 
  x"00",   x"F0",   x"23",   x"D3",   x"46",   x"B6",   x"65",   x"95", 
  x"8C",   x"7C",   x"AF",   x"5F",   x"CA",   x"3A",   x"E9",   x"19", 
  x"DB",   x"2B",   x"F8",   x"08",   x"9D",   x"6D",   x"BE",   x"4E", 
  x"57",   x"A7",   x"74",   x"84",   x"11",   x"E1",   x"32",   x"C2", 
  x"75",   x"85",   x"56",   x"A6",   x"33",   x"C3",   x"10",   x"E0", 
  x"F9",   x"09",   x"DA",   x"2A",   x"BF",   x"4F",   x"9C",   x"6C", 
  x"AE",   x"5E",   x"8D",   x"7D",   x"E8",   x"18",   x"CB",   x"3B", 
  x"22",   x"D2",   x"01",   x"F1",   x"64",   x"94",   x"47",   x"B7", 
  x"EA",   x"1A",   x"C9",   x"39",   x"AC",   x"5C",   x"8F",   x"7F", 
  x"66",   x"96",   x"45",   x"B5",   x"20",   x"D0",   x"03",   x"F3", 
  x"31",   x"C1",   x"12",   x"E2",   x"77",   x"87",   x"54",   x"A4", 
  x"BD",   x"4D",   x"9E",   x"6E",   x"FB",   x"0B",   x"D8",   x"28", 
  x"9F",   x"6F",   x"BC",   x"4C",   x"D9",   x"29",   x"FA",   x"0A", 
  x"13",   x"E3",   x"30",   x"C0",   x"55",   x"A5",   x"76",   x"86", 
  x"44",   x"B4",   x"67",   x"97",   x"02",   x"F2",   x"21",   x"D1", 
  x"C8",   x"38",   x"EB",   x"1B",   x"8E",   x"7E",   x"AD",   x"5D", 
  x"17",   x"E7",   x"34",   x"C4",   x"51",   x"A1",   x"72",   x"82", 
  x"9B",   x"6B",   x"B8",   x"48",   x"DD",   x"2D",   x"FE",   x"0E", 
  x"CC",   x"3C",   x"EF",   x"1F",   x"8A",   x"7A",   x"A9",   x"59", 
  x"40",   x"B0",   x"63",   x"93",   x"06",   x"F6",   x"25",   x"D5", 
  x"62",   x"92",   x"41",   x"B1",   x"24",   x"D4",   x"07",   x"F7", 
  x"EE",   x"1E",   x"CD",   x"3D",   x"A8",   x"58",   x"8B",   x"7B", 
  x"B9",   x"49",   x"9A",   x"6A",   x"FF",   x"0F",   x"DC",   x"2C", 
  x"35",   x"C5",   x"16",   x"E6",   x"73",   x"83",   x"50",   x"A0", 
  x"FD",   x"0D",   x"DE",   x"2E",   x"BB",   x"4B",   x"98",   x"68", 
  x"71",   x"81",   x"52",   x"A2",   x"37",   x"C7",   x"14",   x"E4", 
  x"26",   x"D6",   x"05",   x"F5",   x"60",   x"90",   x"43",   x"B3", 
  x"AA",   x"5A",   x"89",   x"79",   x"EC",   x"1C",   x"CF",   x"3F", 
  x"88",   x"78",   x"AB",   x"5B",   x"CE",   x"3E",   x"ED",   x"1D", 
  x"04",   x"F4",   x"27",   x"D7",   x"42",   x"B2",   x"61",   x"91", 
  x"53",   x"A3",   x"70",   x"80",   x"15",   x"E5",   x"36",   x"C6", 
  x"DF",   x"2F",   x"FC",   x"0C",   x"99",   x"69",   x"BA",   x"4A", 
  x"00",   x"F1",   x"21",   x"D0",   x"42",   x"B3",   x"63",   x"92", 
  x"84",   x"75",   x"A5",   x"54",   x"C6",   x"37",   x"E7",   x"16", 
  x"CB",   x"3A",   x"EA",   x"1B",   x"89",   x"78",   x"A8",   x"59", 
  x"4F",   x"BE",   x"6E",   x"9F",   x"0D",   x"FC",   x"2C",   x"DD", 
  x"55",   x"A4",   x"74",   x"85",   x"17",   x"E6",   x"36",   x"C7", 
  x"D1",   x"20",   x"F0",   x"01",   x"93",   x"62",   x"B2",   x"43", 
  x"9E",   x"6F",   x"BF",   x"4E",   x"DC",   x"2D",   x"FD",   x"0C", 
  x"1A",   x"EB",   x"3B",   x"CA",   x"58",   x"A9",   x"79",   x"88", 
  x"AA",   x"5B",   x"8B",   x"7A",   x"E8",   x"19",   x"C9",   x"38", 
  x"2E",   x"DF",   x"0F",   x"FE",   x"6C",   x"9D",   x"4D",   x"BC", 
  x"61",   x"90",   x"40",   x"B1",   x"23",   x"D2",   x"02",   x"F3", 
  x"E5",   x"14",   x"C4",   x"35",   x"A7",   x"56",   x"86",   x"77", 
  x"FF",   x"0E",   x"DE",   x"2F",   x"BD",   x"4C",   x"9C",   x"6D", 
  x"7B",   x"8A",   x"5A",   x"AB",   x"39",   x"C8",   x"18",   x"E9", 
  x"34",   x"C5",   x"15",   x"E4",   x"76",   x"87",   x"57",   x"A6", 
  x"B0",   x"41",   x"91",   x"60",   x"F2",   x"03",   x"D3",   x"22", 
  x"97",   x"66",   x"B6",   x"47",   x"D5",   x"24",   x"F4",   x"05", 
  x"13",   x"E2",   x"32",   x"C3",   x"51",   x"A0",   x"70",   x"81", 
  x"5C",   x"AD",   x"7D",   x"8C",   x"1E",   x"EF",   x"3F",   x"CE", 
  x"D8",   x"29",   x"F9",   x"08",   x"9A",   x"6B",   x"BB",   x"4A", 
  x"C2",   x"33",   x"E3",   x"12",   x"80",   x"71",   x"A1",   x"50", 
  x"46",   x"B7",   x"67",   x"96",   x"04",   x"F5",   x"25",   x"D4", 
  x"09",   x"F8",   x"28",   x"D9",   x"4B",   x"BA",   x"6A",   x"9B", 
  x"8D",   x"7C",   x"AC",   x"5D",   x"CF",   x"3E",   x"EE",   x"1F", 
  x"3D",   x"CC",   x"1C",   x"ED",   x"7F",   x"8E",   x"5E",   x"AF", 
  x"B9",   x"48",   x"98",   x"69",   x"FB",   x"0A",   x"DA",   x"2B", 
  x"F6",   x"07",   x"D7",   x"26",   x"B4",   x"45",   x"95",   x"64", 
  x"72",   x"83",   x"53",   x"A2",   x"30",   x"C1",   x"11",   x"E0", 
  x"68",   x"99",   x"49",   x"B8",   x"2A",   x"DB",   x"0B",   x"FA", 
  x"EC",   x"1D",   x"CD",   x"3C",   x"AE",   x"5F",   x"8F",   x"7E", 
  x"A3",   x"52",   x"82",   x"73",   x"E1",   x"10",   x"C0",   x"31", 
  x"27",   x"D6",   x"06",   x"F7",   x"65",   x"94",   x"44",   x"B5", 
  x"00",   x"F2",   x"27",   x"D5",   x"4E",   x"BC",   x"69",   x"9B", 
  x"9C",   x"6E",   x"BB",   x"49",   x"D2",   x"20",   x"F5",   x"07", 
  x"FB",   x"09",   x"DC",   x"2E",   x"B5",   x"47",   x"92",   x"60", 
  x"67",   x"95",   x"40",   x"B2",   x"29",   x"DB",   x"0E",   x"FC", 
  x"35",   x"C7",   x"12",   x"E0",   x"7B",   x"89",   x"5C",   x"AE", 
  x"A9",   x"5B",   x"8E",   x"7C",   x"E7",   x"15",   x"C0",   x"32", 
  x"CE",   x"3C",   x"E9",   x"1B",   x"80",   x"72",   x"A7",   x"55", 
  x"52",   x"A0",   x"75",   x"87",   x"1C",   x"EE",   x"3B",   x"C9", 
  x"6A",   x"98",   x"4D",   x"BF",   x"24",   x"D6",   x"03",   x"F1", 
  x"F6",   x"04",   x"D1",   x"23",   x"B8",   x"4A",   x"9F",   x"6D", 
  x"91",   x"63",   x"B6",   x"44",   x"DF",   x"2D",   x"F8",   x"0A", 
  x"0D",   x"FF",   x"2A",   x"D8",   x"43",   x"B1",   x"64",   x"96", 
  x"5F",   x"AD",   x"78",   x"8A",   x"11",   x"E3",   x"36",   x"C4", 
  x"C3",   x"31",   x"E4",   x"16",   x"8D",   x"7F",   x"AA",   x"58", 
  x"A4",   x"56",   x"83",   x"71",   x"EA",   x"18",   x"CD",   x"3F", 
  x"38",   x"CA",   x"1F",   x"ED",   x"76",   x"84",   x"51",   x"A3", 
  x"D4",   x"26",   x"F3",   x"01",   x"9A",   x"68",   x"BD",   x"4F", 
  x"48",   x"BA",   x"6F",   x"9D",   x"06",   x"F4",   x"21",   x"D3", 
  x"2F",   x"DD",   x"08",   x"FA",   x"61",   x"93",   x"46",   x"B4", 
  x"B3",   x"41",   x"94",   x"66",   x"FD",   x"0F",   x"DA",   x"28", 
  x"E1",   x"13",   x"C6",   x"34",   x"AF",   x"5D",   x"88",   x"7A", 
  x"7D",   x"8F",   x"5A",   x"A8",   x"33",   x"C1",   x"14",   x"E6", 
  x"1A",   x"E8",   x"3D",   x"CF",   x"54",   x"A6",   x"73",   x"81", 
  x"86",   x"74",   x"A1",   x"53",   x"C8",   x"3A",   x"EF",   x"1D", 
  x"BE",   x"4C",   x"99",   x"6B",   x"F0",   x"02",   x"D7",   x"25", 
  x"22",   x"D0",   x"05",   x"F7",   x"6C",   x"9E",   x"4B",   x"B9", 
  x"45",   x"B7",   x"62",   x"90",   x"0B",   x"F9",   x"2C",   x"DE", 
  x"D9",   x"2B",   x"FE",   x"0C",   x"97",   x"65",   x"B0",   x"42", 
  x"8B",   x"79",   x"AC",   x"5E",   x"C5",   x"37",   x"E2",   x"10", 
  x"17",   x"E5",   x"30",   x"C2",   x"59",   x"AB",   x"7E",   x"8C", 
  x"70",   x"82",   x"57",   x"A5",   x"3E",   x"CC",   x"19",   x"EB", 
  x"EC",   x"1E",   x"CB",   x"39",   x"A2",   x"50",   x"85",   x"77", 
  x"00",   x"F3",   x"25",   x"D6",   x"4A",   x"B9",   x"6F",   x"9C", 
  x"94",   x"67",   x"B1",   x"42",   x"DE",   x"2D",   x"FB",   x"08", 
  x"EB",   x"18",   x"CE",   x"3D",   x"A1",   x"52",   x"84",   x"77", 
  x"7F",   x"8C",   x"5A",   x"A9",   x"35",   x"C6",   x"10",   x"E3", 
  x"15",   x"E6",   x"30",   x"C3",   x"5F",   x"AC",   x"7A",   x"89", 
  x"81",   x"72",   x"A4",   x"57",   x"CB",   x"38",   x"EE",   x"1D", 
  x"FE",   x"0D",   x"DB",   x"28",   x"B4",   x"47",   x"91",   x"62", 
  x"6A",   x"99",   x"4F",   x"BC",   x"20",   x"D3",   x"05",   x"F6", 
  x"2A",   x"D9",   x"0F",   x"FC",   x"60",   x"93",   x"45",   x"B6", 
  x"BE",   x"4D",   x"9B",   x"68",   x"F4",   x"07",   x"D1",   x"22", 
  x"C1",   x"32",   x"E4",   x"17",   x"8B",   x"78",   x"AE",   x"5D", 
  x"55",   x"A6",   x"70",   x"83",   x"1F",   x"EC",   x"3A",   x"C9", 
  x"3F",   x"CC",   x"1A",   x"E9",   x"75",   x"86",   x"50",   x"A3", 
  x"AB",   x"58",   x"8E",   x"7D",   x"E1",   x"12",   x"C4",   x"37", 
  x"D4",   x"27",   x"F1",   x"02",   x"9E",   x"6D",   x"BB",   x"48", 
  x"40",   x"B3",   x"65",   x"96",   x"0A",   x"F9",   x"2F",   x"DC", 
  x"54",   x"A7",   x"71",   x"82",   x"1E",   x"ED",   x"3B",   x"C8", 
  x"C0",   x"33",   x"E5",   x"16",   x"8A",   x"79",   x"AF",   x"5C", 
  x"BF",   x"4C",   x"9A",   x"69",   x"F5",   x"06",   x"D0",   x"23", 
  x"2B",   x"D8",   x"0E",   x"FD",   x"61",   x"92",   x"44",   x"B7", 
  x"41",   x"B2",   x"64",   x"97",   x"0B",   x"F8",   x"2E",   x"DD", 
  x"D5",   x"26",   x"F0",   x"03",   x"9F",   x"6C",   x"BA",   x"49", 
  x"AA",   x"59",   x"8F",   x"7C",   x"E0",   x"13",   x"C5",   x"36", 
  x"3E",   x"CD",   x"1B",   x"E8",   x"74",   x"87",   x"51",   x"A2", 
  x"7E",   x"8D",   x"5B",   x"A8",   x"34",   x"C7",   x"11",   x"E2", 
  x"EA",   x"19",   x"CF",   x"3C",   x"A0",   x"53",   x"85",   x"76", 
  x"95",   x"66",   x"B0",   x"43",   x"DF",   x"2C",   x"FA",   x"09", 
  x"01",   x"F2",   x"24",   x"D7",   x"4B",   x"B8",   x"6E",   x"9D", 
  x"6B",   x"98",   x"4E",   x"BD",   x"21",   x"D2",   x"04",   x"F7", 
  x"FF",   x"0C",   x"DA",   x"29",   x"B5",   x"46",   x"90",   x"63", 
  x"80",   x"73",   x"A5",   x"56",   x"CA",   x"39",   x"EF",   x"1C", 
  x"14",   x"E7",   x"31",   x"C2",   x"5E",   x"AD",   x"7B",   x"88", 
  x"00",   x"F4",   x"2B",   x"DF",   x"56",   x"A2",   x"7D",   x"89", 
  x"AC",   x"58",   x"87",   x"73",   x"FA",   x"0E",   x"D1",   x"25", 
  x"9B",   x"6F",   x"B0",   x"44",   x"CD",   x"39",   x"E6",   x"12", 
  x"37",   x"C3",   x"1C",   x"E8",   x"61",   x"95",   x"4A",   x"BE", 
  x"F5",   x"01",   x"DE",   x"2A",   x"A3",   x"57",   x"88",   x"7C", 
  x"59",   x"AD",   x"72",   x"86",   x"0F",   x"FB",   x"24",   x"D0", 
  x"6E",   x"9A",   x"45",   x"B1",   x"38",   x"CC",   x"13",   x"E7", 
  x"C2",   x"36",   x"E9",   x"1D",   x"94",   x"60",   x"BF",   x"4B", 
  x"29",   x"DD",   x"02",   x"F6",   x"7F",   x"8B",   x"54",   x"A0", 
  x"85",   x"71",   x"AE",   x"5A",   x"D3",   x"27",   x"F8",   x"0C", 
  x"B2",   x"46",   x"99",   x"6D",   x"E4",   x"10",   x"CF",   x"3B", 
  x"1E",   x"EA",   x"35",   x"C1",   x"48",   x"BC",   x"63",   x"97", 
  x"DC",   x"28",   x"F7",   x"03",   x"8A",   x"7E",   x"A1",   x"55", 
  x"70",   x"84",   x"5B",   x"AF",   x"26",   x"D2",   x"0D",   x"F9", 
  x"47",   x"B3",   x"6C",   x"98",   x"11",   x"E5",   x"3A",   x"CE", 
  x"EB",   x"1F",   x"C0",   x"34",   x"BD",   x"49",   x"96",   x"62", 
  x"52",   x"A6",   x"79",   x"8D",   x"04",   x"F0",   x"2F",   x"DB", 
  x"FE",   x"0A",   x"D5",   x"21",   x"A8",   x"5C",   x"83",   x"77", 
  x"C9",   x"3D",   x"E2",   x"16",   x"9F",   x"6B",   x"B4",   x"40", 
  x"65",   x"91",   x"4E",   x"BA",   x"33",   x"C7",   x"18",   x"EC", 
  x"A7",   x"53",   x"8C",   x"78",   x"F1",   x"05",   x"DA",   x"2E", 
  x"0B",   x"FF",   x"20",   x"D4",   x"5D",   x"A9",   x"76",   x"82", 
  x"3C",   x"C8",   x"17",   x"E3",   x"6A",   x"9E",   x"41",   x"B5", 
  x"90",   x"64",   x"BB",   x"4F",   x"C6",   x"32",   x"ED",   x"19", 
  x"7B",   x"8F",   x"50",   x"A4",   x"2D",   x"D9",   x"06",   x"F2", 
  x"D7",   x"23",   x"FC",   x"08",   x"81",   x"75",   x"AA",   x"5E", 
  x"E0",   x"14",   x"CB",   x"3F",   x"B6",   x"42",   x"9D",   x"69", 
  x"4C",   x"B8",   x"67",   x"93",   x"1A",   x"EE",   x"31",   x"C5", 
  x"8E",   x"7A",   x"A5",   x"51",   x"D8",   x"2C",   x"F3",   x"07", 
  x"22",   x"D6",   x"09",   x"FD",   x"74",   x"80",   x"5F",   x"AB", 
  x"15",   x"E1",   x"3E",   x"CA",   x"43",   x"B7",   x"68",   x"9C", 
  x"B9",   x"4D",   x"92",   x"66",   x"EF",   x"1B",   x"C4",   x"30", 
  x"00",   x"F5",   x"29",   x"DC",   x"52",   x"A7",   x"7B",   x"8E", 
  x"A4",   x"51",   x"8D",   x"78",   x"F6",   x"03",   x"DF",   x"2A", 
  x"8B",   x"7E",   x"A2",   x"57",   x"D9",   x"2C",   x"F0",   x"05", 
  x"2F",   x"DA",   x"06",   x"F3",   x"7D",   x"88",   x"54",   x"A1", 
  x"D5",   x"20",   x"FC",   x"09",   x"87",   x"72",   x"AE",   x"5B", 
  x"71",   x"84",   x"58",   x"AD",   x"23",   x"D6",   x"0A",   x"FF", 
  x"5E",   x"AB",   x"77",   x"82",   x"0C",   x"F9",   x"25",   x"D0", 
  x"FA",   x"0F",   x"D3",   x"26",   x"A8",   x"5D",   x"81",   x"74", 
  x"69",   x"9C",   x"40",   x"B5",   x"3B",   x"CE",   x"12",   x"E7", 
  x"CD",   x"38",   x"E4",   x"11",   x"9F",   x"6A",   x"B6",   x"43", 
  x"E2",   x"17",   x"CB",   x"3E",   x"B0",   x"45",   x"99",   x"6C", 
  x"46",   x"B3",   x"6F",   x"9A",   x"14",   x"E1",   x"3D",   x"C8", 
  x"BC",   x"49",   x"95",   x"60",   x"EE",   x"1B",   x"C7",   x"32", 
  x"18",   x"ED",   x"31",   x"C4",   x"4A",   x"BF",   x"63",   x"96", 
  x"37",   x"C2",   x"1E",   x"EB",   x"65",   x"90",   x"4C",   x"B9", 
  x"93",   x"66",   x"BA",   x"4F",   x"C1",   x"34",   x"E8",   x"1D", 
  x"D2",   x"27",   x"FB",   x"0E",   x"80",   x"75",   x"A9",   x"5C", 
  x"76",   x"83",   x"5F",   x"AA",   x"24",   x"D1",   x"0D",   x"F8", 
  x"59",   x"AC",   x"70",   x"85",   x"0B",   x"FE",   x"22",   x"D7", 
  x"FD",   x"08",   x"D4",   x"21",   x"AF",   x"5A",   x"86",   x"73", 
  x"07",   x"F2",   x"2E",   x"DB",   x"55",   x"A0",   x"7C",   x"89", 
  x"A3",   x"56",   x"8A",   x"7F",   x"F1",   x"04",   x"D8",   x"2D", 
  x"8C",   x"79",   x"A5",   x"50",   x"DE",   x"2B",   x"F7",   x"02", 
  x"28",   x"DD",   x"01",   x"F4",   x"7A",   x"8F",   x"53",   x"A6", 
  x"BB",   x"4E",   x"92",   x"67",   x"E9",   x"1C",   x"C0",   x"35", 
  x"1F",   x"EA",   x"36",   x"C3",   x"4D",   x"B8",   x"64",   x"91", 
  x"30",   x"C5",   x"19",   x"EC",   x"62",   x"97",   x"4B",   x"BE", 
  x"94",   x"61",   x"BD",   x"48",   x"C6",   x"33",   x"EF",   x"1A", 
  x"6E",   x"9B",   x"47",   x"B2",   x"3C",   x"C9",   x"15",   x"E0", 
  x"CA",   x"3F",   x"E3",   x"16",   x"98",   x"6D",   x"B1",   x"44", 
  x"E5",   x"10",   x"CC",   x"39",   x"B7",   x"42",   x"9E",   x"6B", 
  x"41",   x"B4",   x"68",   x"9D",   x"13",   x"E6",   x"3A",   x"CF", 
  x"00",   x"F6",   x"2F",   x"D9",   x"5E",   x"A8",   x"71",   x"87", 
  x"BC",   x"4A",   x"93",   x"65",   x"E2",   x"14",   x"CD",   x"3B", 
  x"BB",   x"4D",   x"94",   x"62",   x"E5",   x"13",   x"CA",   x"3C", 
  x"07",   x"F1",   x"28",   x"DE",   x"59",   x"AF",   x"76",   x"80", 
  x"B5",   x"43",   x"9A",   x"6C",   x"EB",   x"1D",   x"C4",   x"32", 
  x"09",   x"FF",   x"26",   x"D0",   x"57",   x"A1",   x"78",   x"8E", 
  x"0E",   x"F8",   x"21",   x"D7",   x"50",   x"A6",   x"7F",   x"89", 
  x"B2",   x"44",   x"9D",   x"6B",   x"EC",   x"1A",   x"C3",   x"35", 
  x"A9",   x"5F",   x"86",   x"70",   x"F7",   x"01",   x"D8",   x"2E", 
  x"15",   x"E3",   x"3A",   x"CC",   x"4B",   x"BD",   x"64",   x"92", 
  x"12",   x"E4",   x"3D",   x"CB",   x"4C",   x"BA",   x"63",   x"95", 
  x"AE",   x"58",   x"81",   x"77",   x"F0",   x"06",   x"DF",   x"29", 
  x"1C",   x"EA",   x"33",   x"C5",   x"42",   x"B4",   x"6D",   x"9B", 
  x"A0",   x"56",   x"8F",   x"79",   x"FE",   x"08",   x"D1",   x"27", 
  x"A7",   x"51",   x"88",   x"7E",   x"F9",   x"0F",   x"D6",   x"20", 
  x"1B",   x"ED",   x"34",   x"C2",   x"45",   x"B3",   x"6A",   x"9C", 
  x"91",   x"67",   x"BE",   x"48",   x"CF",   x"39",   x"E0",   x"16", 
  x"2D",   x"DB",   x"02",   x"F4",   x"73",   x"85",   x"5C",   x"AA", 
  x"2A",   x"DC",   x"05",   x"F3",   x"74",   x"82",   x"5B",   x"AD", 
  x"96",   x"60",   x"B9",   x"4F",   x"C8",   x"3E",   x"E7",   x"11", 
  x"24",   x"D2",   x"0B",   x"FD",   x"7A",   x"8C",   x"55",   x"A3", 
  x"98",   x"6E",   x"B7",   x"41",   x"C6",   x"30",   x"E9",   x"1F", 
  x"9F",   x"69",   x"B0",   x"46",   x"C1",   x"37",   x"EE",   x"18", 
  x"23",   x"D5",   x"0C",   x"FA",   x"7D",   x"8B",   x"52",   x"A4", 
  x"38",   x"CE",   x"17",   x"E1",   x"66",   x"90",   x"49",   x"BF", 
  x"84",   x"72",   x"AB",   x"5D",   x"DA",   x"2C",   x"F5",   x"03", 
  x"83",   x"75",   x"AC",   x"5A",   x"DD",   x"2B",   x"F2",   x"04", 
  x"3F",   x"C9",   x"10",   x"E6",   x"61",   x"97",   x"4E",   x"B8", 
  x"8D",   x"7B",   x"A2",   x"54",   x"D3",   x"25",   x"FC",   x"0A", 
  x"31",   x"C7",   x"1E",   x"E8",   x"6F",   x"99",   x"40",   x"B6", 
  x"36",   x"C0",   x"19",   x"EF",   x"68",   x"9E",   x"47",   x"B1", 
  x"8A",   x"7C",   x"A5",   x"53",   x"D4",   x"22",   x"FB",   x"0D", 
  x"00",   x"F7",   x"2D",   x"DA",   x"5A",   x"AD",   x"77",   x"80", 
  x"B4",   x"43",   x"99",   x"6E",   x"EE",   x"19",   x"C3",   x"34", 
  x"AB",   x"5C",   x"86",   x"71",   x"F1",   x"06",   x"DC",   x"2B", 
  x"1F",   x"E8",   x"32",   x"C5",   x"45",   x"B2",   x"68",   x"9F", 
  x"95",   x"62",   x"B8",   x"4F",   x"CF",   x"38",   x"E2",   x"15", 
  x"21",   x"D6",   x"0C",   x"FB",   x"7B",   x"8C",   x"56",   x"A1", 
  x"3E",   x"C9",   x"13",   x"E4",   x"64",   x"93",   x"49",   x"BE", 
  x"8A",   x"7D",   x"A7",   x"50",   x"D0",   x"27",   x"FD",   x"0A", 
  x"E9",   x"1E",   x"C4",   x"33",   x"B3",   x"44",   x"9E",   x"69", 
  x"5D",   x"AA",   x"70",   x"87",   x"07",   x"F0",   x"2A",   x"DD", 
  x"42",   x"B5",   x"6F",   x"98",   x"18",   x"EF",   x"35",   x"C2", 
  x"F6",   x"01",   x"DB",   x"2C",   x"AC",   x"5B",   x"81",   x"76", 
  x"7C",   x"8B",   x"51",   x"A6",   x"26",   x"D1",   x"0B",   x"FC", 
  x"C8",   x"3F",   x"E5",   x"12",   x"92",   x"65",   x"BF",   x"48", 
  x"D7",   x"20",   x"FA",   x"0D",   x"8D",   x"7A",   x"A0",   x"57", 
  x"63",   x"94",   x"4E",   x"B9",   x"39",   x"CE",   x"14",   x"E3", 
  x"11",   x"E6",   x"3C",   x"CB",   x"4B",   x"BC",   x"66",   x"91", 
  x"A5",   x"52",   x"88",   x"7F",   x"FF",   x"08",   x"D2",   x"25", 
  x"BA",   x"4D",   x"97",   x"60",   x"E0",   x"17",   x"CD",   x"3A", 
  x"0E",   x"F9",   x"23",   x"D4",   x"54",   x"A3",   x"79",   x"8E", 
  x"84",   x"73",   x"A9",   x"5E",   x"DE",   x"29",   x"F3",   x"04", 
  x"30",   x"C7",   x"1D",   x"EA",   x"6A",   x"9D",   x"47",   x"B0", 
  x"2F",   x"D8",   x"02",   x"F5",   x"75",   x"82",   x"58",   x"AF", 
  x"9B",   x"6C",   x"B6",   x"41",   x"C1",   x"36",   x"EC",   x"1B", 
  x"F8",   x"0F",   x"D5",   x"22",   x"A2",   x"55",   x"8F",   x"78", 
  x"4C",   x"BB",   x"61",   x"96",   x"16",   x"E1",   x"3B",   x"CC", 
  x"53",   x"A4",   x"7E",   x"89",   x"09",   x"FE",   x"24",   x"D3", 
  x"E7",   x"10",   x"CA",   x"3D",   x"BD",   x"4A",   x"90",   x"67", 
  x"6D",   x"9A",   x"40",   x"B7",   x"37",   x"C0",   x"1A",   x"ED", 
  x"D9",   x"2E",   x"F4",   x"03",   x"83",   x"74",   x"AE",   x"59", 
  x"C6",   x"31",   x"EB",   x"1C",   x"9C",   x"6B",   x"B1",   x"46", 
  x"72",   x"85",   x"5F",   x"A8",   x"28",   x"DF",   x"05",   x"F2", 
  x"00",   x"F8",   x"33",   x"CB",   x"66",   x"9E",   x"55",   x"AD", 
  x"CC",   x"34",   x"FF",   x"07",   x"AA",   x"52",   x"99",   x"61", 
  x"5B",   x"A3",   x"68",   x"90",   x"3D",   x"C5",   x"0E",   x"F6", 
  x"97",   x"6F",   x"A4",   x"5C",   x"F1",   x"09",   x"C2",   x"3A", 
  x"B6",   x"4E",   x"85",   x"7D",   x"D0",   x"28",   x"E3",   x"1B", 
  x"7A",   x"82",   x"49",   x"B1",   x"1C",   x"E4",   x"2F",   x"D7", 
  x"ED",   x"15",   x"DE",   x"26",   x"8B",   x"73",   x"B8",   x"40", 
  x"21",   x"D9",   x"12",   x"EA",   x"47",   x"BF",   x"74",   x"8C", 
  x"AF",   x"57",   x"9C",   x"64",   x"C9",   x"31",   x"FA",   x"02", 
  x"63",   x"9B",   x"50",   x"A8",   x"05",   x"FD",   x"36",   x"CE", 
  x"F4",   x"0C",   x"C7",   x"3F",   x"92",   x"6A",   x"A1",   x"59", 
  x"38",   x"C0",   x"0B",   x"F3",   x"5E",   x"A6",   x"6D",   x"95", 
  x"19",   x"E1",   x"2A",   x"D2",   x"7F",   x"87",   x"4C",   x"B4", 
  x"D5",   x"2D",   x"E6",   x"1E",   x"B3",   x"4B",   x"80",   x"78", 
  x"42",   x"BA",   x"71",   x"89",   x"24",   x"DC",   x"17",   x"EF", 
  x"8E",   x"76",   x"BD",   x"45",   x"E8",   x"10",   x"DB",   x"23", 
  x"9D",   x"65",   x"AE",   x"56",   x"FB",   x"03",   x"C8",   x"30", 
  x"51",   x"A9",   x"62",   x"9A",   x"37",   x"CF",   x"04",   x"FC", 
  x"C6",   x"3E",   x"F5",   x"0D",   x"A0",   x"58",   x"93",   x"6B", 
  x"0A",   x"F2",   x"39",   x"C1",   x"6C",   x"94",   x"5F",   x"A7", 
  x"2B",   x"D3",   x"18",   x"E0",   x"4D",   x"B5",   x"7E",   x"86", 
  x"E7",   x"1F",   x"D4",   x"2C",   x"81",   x"79",   x"B2",   x"4A", 
  x"70",   x"88",   x"43",   x"BB",   x"16",   x"EE",   x"25",   x"DD", 
  x"BC",   x"44",   x"8F",   x"77",   x"DA",   x"22",   x"E9",   x"11", 
  x"32",   x"CA",   x"01",   x"F9",   x"54",   x"AC",   x"67",   x"9F", 
  x"FE",   x"06",   x"CD",   x"35",   x"98",   x"60",   x"AB",   x"53", 
  x"69",   x"91",   x"5A",   x"A2",   x"0F",   x"F7",   x"3C",   x"C4", 
  x"A5",   x"5D",   x"96",   x"6E",   x"C3",   x"3B",   x"F0",   x"08", 
  x"84",   x"7C",   x"B7",   x"4F",   x"E2",   x"1A",   x"D1",   x"29", 
  x"48",   x"B0",   x"7B",   x"83",   x"2E",   x"D6",   x"1D",   x"E5", 
  x"DF",   x"27",   x"EC",   x"14",   x"B9",   x"41",   x"8A",   x"72", 
  x"13",   x"EB",   x"20",   x"D8",   x"75",   x"8D",   x"46",   x"BE", 
  x"00",   x"F9",   x"31",   x"C8",   x"62",   x"9B",   x"53",   x"AA", 
  x"C4",   x"3D",   x"F5",   x"0C",   x"A6",   x"5F",   x"97",   x"6E", 
  x"4B",   x"B2",   x"7A",   x"83",   x"29",   x"D0",   x"18",   x"E1", 
  x"8F",   x"76",   x"BE",   x"47",   x"ED",   x"14",   x"DC",   x"25", 
  x"96",   x"6F",   x"A7",   x"5E",   x"F4",   x"0D",   x"C5",   x"3C", 
  x"52",   x"AB",   x"63",   x"9A",   x"30",   x"C9",   x"01",   x"F8", 
  x"DD",   x"24",   x"EC",   x"15",   x"BF",   x"46",   x"8E",   x"77", 
  x"19",   x"E0",   x"28",   x"D1",   x"7B",   x"82",   x"4A",   x"B3", 
  x"EF",   x"16",   x"DE",   x"27",   x"8D",   x"74",   x"BC",   x"45", 
  x"2B",   x"D2",   x"1A",   x"E3",   x"49",   x"B0",   x"78",   x"81", 
  x"A4",   x"5D",   x"95",   x"6C",   x"C6",   x"3F",   x"F7",   x"0E", 
  x"60",   x"99",   x"51",   x"A8",   x"02",   x"FB",   x"33",   x"CA", 
  x"79",   x"80",   x"48",   x"B1",   x"1B",   x"E2",   x"2A",   x"D3", 
  x"BD",   x"44",   x"8C",   x"75",   x"DF",   x"26",   x"EE",   x"17", 
  x"32",   x"CB",   x"03",   x"FA",   x"50",   x"A9",   x"61",   x"98", 
  x"F6",   x"0F",   x"C7",   x"3E",   x"94",   x"6D",   x"A5",   x"5C", 
  x"1D",   x"E4",   x"2C",   x"D5",   x"7F",   x"86",   x"4E",   x"B7", 
  x"D9",   x"20",   x"E8",   x"11",   x"BB",   x"42",   x"8A",   x"73", 
  x"56",   x"AF",   x"67",   x"9E",   x"34",   x"CD",   x"05",   x"FC", 
  x"92",   x"6B",   x"A3",   x"5A",   x"F0",   x"09",   x"C1",   x"38", 
  x"8B",   x"72",   x"BA",   x"43",   x"E9",   x"10",   x"D8",   x"21", 
  x"4F",   x"B6",   x"7E",   x"87",   x"2D",   x"D4",   x"1C",   x"E5", 
  x"C0",   x"39",   x"F1",   x"08",   x"A2",   x"5B",   x"93",   x"6A", 
  x"04",   x"FD",   x"35",   x"CC",   x"66",   x"9F",   x"57",   x"AE", 
  x"F2",   x"0B",   x"C3",   x"3A",   x"90",   x"69",   x"A1",   x"58", 
  x"36",   x"CF",   x"07",   x"FE",   x"54",   x"AD",   x"65",   x"9C", 
  x"B9",   x"40",   x"88",   x"71",   x"DB",   x"22",   x"EA",   x"13", 
  x"7D",   x"84",   x"4C",   x"B5",   x"1F",   x"E6",   x"2E",   x"D7", 
  x"64",   x"9D",   x"55",   x"AC",   x"06",   x"FF",   x"37",   x"CE", 
  x"A0",   x"59",   x"91",   x"68",   x"C2",   x"3B",   x"F3",   x"0A", 
  x"2F",   x"D6",   x"1E",   x"E7",   x"4D",   x"B4",   x"7C",   x"85", 
  x"EB",   x"12",   x"DA",   x"23",   x"89",   x"70",   x"B8",   x"41", 
  x"00",   x"FA",   x"37",   x"CD",   x"6E",   x"94",   x"59",   x"A3", 
  x"DC",   x"26",   x"EB",   x"11",   x"B2",   x"48",   x"85",   x"7F", 
  x"7B",   x"81",   x"4C",   x"B6",   x"15",   x"EF",   x"22",   x"D8", 
  x"A7",   x"5D",   x"90",   x"6A",   x"C9",   x"33",   x"FE",   x"04", 
  x"F6",   x"0C",   x"C1",   x"3B",   x"98",   x"62",   x"AF",   x"55", 
  x"2A",   x"D0",   x"1D",   x"E7",   x"44",   x"BE",   x"73",   x"89", 
  x"8D",   x"77",   x"BA",   x"40",   x"E3",   x"19",   x"D4",   x"2E", 
  x"51",   x"AB",   x"66",   x"9C",   x"3F",   x"C5",   x"08",   x"F2", 
  x"2F",   x"D5",   x"18",   x"E2",   x"41",   x"BB",   x"76",   x"8C", 
  x"F3",   x"09",   x"C4",   x"3E",   x"9D",   x"67",   x"AA",   x"50", 
  x"54",   x"AE",   x"63",   x"99",   x"3A",   x"C0",   x"0D",   x"F7", 
  x"88",   x"72",   x"BF",   x"45",   x"E6",   x"1C",   x"D1",   x"2B", 
  x"D9",   x"23",   x"EE",   x"14",   x"B7",   x"4D",   x"80",   x"7A", 
  x"05",   x"FF",   x"32",   x"C8",   x"6B",   x"91",   x"5C",   x"A6", 
  x"A2",   x"58",   x"95",   x"6F",   x"CC",   x"36",   x"FB",   x"01", 
  x"7E",   x"84",   x"49",   x"B3",   x"10",   x"EA",   x"27",   x"DD", 
  x"5E",   x"A4",   x"69",   x"93",   x"30",   x"CA",   x"07",   x"FD", 
  x"82",   x"78",   x"B5",   x"4F",   x"EC",   x"16",   x"DB",   x"21", 
  x"25",   x"DF",   x"12",   x"E8",   x"4B",   x"B1",   x"7C",   x"86", 
  x"F9",   x"03",   x"CE",   x"34",   x"97",   x"6D",   x"A0",   x"5A", 
  x"A8",   x"52",   x"9F",   x"65",   x"C6",   x"3C",   x"F1",   x"0B", 
  x"74",   x"8E",   x"43",   x"B9",   x"1A",   x"E0",   x"2D",   x"D7", 
  x"D3",   x"29",   x"E4",   x"1E",   x"BD",   x"47",   x"8A",   x"70", 
  x"0F",   x"F5",   x"38",   x"C2",   x"61",   x"9B",   x"56",   x"AC", 
  x"71",   x"8B",   x"46",   x"BC",   x"1F",   x"E5",   x"28",   x"D2", 
  x"AD",   x"57",   x"9A",   x"60",   x"C3",   x"39",   x"F4",   x"0E", 
  x"0A",   x"F0",   x"3D",   x"C7",   x"64",   x"9E",   x"53",   x"A9", 
  x"D6",   x"2C",   x"E1",   x"1B",   x"B8",   x"42",   x"8F",   x"75", 
  x"87",   x"7D",   x"B0",   x"4A",   x"E9",   x"13",   x"DE",   x"24", 
  x"5B",   x"A1",   x"6C",   x"96",   x"35",   x"CF",   x"02",   x"F8", 
  x"FC",   x"06",   x"CB",   x"31",   x"92",   x"68",   x"A5",   x"5F", 
  x"20",   x"DA",   x"17",   x"ED",   x"4E",   x"B4",   x"79",   x"83", 
  x"00",   x"FB",   x"35",   x"CE",   x"6A",   x"91",   x"5F",   x"A4", 
  x"D4",   x"2F",   x"E1",   x"1A",   x"BE",   x"45",   x"8B",   x"70", 
  x"6B",   x"90",   x"5E",   x"A5",   x"01",   x"FA",   x"34",   x"CF", 
  x"BF",   x"44",   x"8A",   x"71",   x"D5",   x"2E",   x"E0",   x"1B", 
  x"D6",   x"2D",   x"E3",   x"18",   x"BC",   x"47",   x"89",   x"72", 
  x"02",   x"F9",   x"37",   x"CC",   x"68",   x"93",   x"5D",   x"A6", 
  x"BD",   x"46",   x"88",   x"73",   x"D7",   x"2C",   x"E2",   x"19", 
  x"69",   x"92",   x"5C",   x"A7",   x"03",   x"F8",   x"36",   x"CD", 
  x"6F",   x"94",   x"5A",   x"A1",   x"05",   x"FE",   x"30",   x"CB", 
  x"BB",   x"40",   x"8E",   x"75",   x"D1",   x"2A",   x"E4",   x"1F", 
  x"04",   x"FF",   x"31",   x"CA",   x"6E",   x"95",   x"5B",   x"A0", 
  x"D0",   x"2B",   x"E5",   x"1E",   x"BA",   x"41",   x"8F",   x"74", 
  x"B9",   x"42",   x"8C",   x"77",   x"D3",   x"28",   x"E6",   x"1D", 
  x"6D",   x"96",   x"58",   x"A3",   x"07",   x"FC",   x"32",   x"C9", 
  x"D2",   x"29",   x"E7",   x"1C",   x"B8",   x"43",   x"8D",   x"76", 
  x"06",   x"FD",   x"33",   x"C8",   x"6C",   x"97",   x"59",   x"A2", 
  x"DE",   x"25",   x"EB",   x"10",   x"B4",   x"4F",   x"81",   x"7A", 
  x"0A",   x"F1",   x"3F",   x"C4",   x"60",   x"9B",   x"55",   x"AE", 
  x"B5",   x"4E",   x"80",   x"7B",   x"DF",   x"24",   x"EA",   x"11", 
  x"61",   x"9A",   x"54",   x"AF",   x"0B",   x"F0",   x"3E",   x"C5", 
  x"08",   x"F3",   x"3D",   x"C6",   x"62",   x"99",   x"57",   x"AC", 
  x"DC",   x"27",   x"E9",   x"12",   x"B6",   x"4D",   x"83",   x"78", 
  x"63",   x"98",   x"56",   x"AD",   x"09",   x"F2",   x"3C",   x"C7", 
  x"B7",   x"4C",   x"82",   x"79",   x"DD",   x"26",   x"E8",   x"13", 
  x"B1",   x"4A",   x"84",   x"7F",   x"DB",   x"20",   x"EE",   x"15", 
  x"65",   x"9E",   x"50",   x"AB",   x"0F",   x"F4",   x"3A",   x"C1", 
  x"DA",   x"21",   x"EF",   x"14",   x"B0",   x"4B",   x"85",   x"7E", 
  x"0E",   x"F5",   x"3B",   x"C0",   x"64",   x"9F",   x"51",   x"AA", 
  x"67",   x"9C",   x"52",   x"A9",   x"0D",   x"F6",   x"38",   x"C3", 
  x"B3",   x"48",   x"86",   x"7D",   x"D9",   x"22",   x"EC",   x"17", 
  x"0C",   x"F7",   x"39",   x"C2",   x"66",   x"9D",   x"53",   x"A8", 
  x"D8",   x"23",   x"ED",   x"16",   x"B2",   x"49",   x"87",   x"7C", 
  x"00",   x"FC",   x"3B",   x"C7",   x"76",   x"8A",   x"4D",   x"B1", 
  x"EC",   x"10",   x"D7",   x"2B",   x"9A",   x"66",   x"A1",   x"5D", 
  x"1B",   x"E7",   x"20",   x"DC",   x"6D",   x"91",   x"56",   x"AA", 
  x"F7",   x"0B",   x"CC",   x"30",   x"81",   x"7D",   x"BA",   x"46", 
  x"36",   x"CA",   x"0D",   x"F1",   x"40",   x"BC",   x"7B",   x"87", 
  x"DA",   x"26",   x"E1",   x"1D",   x"AC",   x"50",   x"97",   x"6B", 
  x"2D",   x"D1",   x"16",   x"EA",   x"5B",   x"A7",   x"60",   x"9C", 
  x"C1",   x"3D",   x"FA",   x"06",   x"B7",   x"4B",   x"8C",   x"70", 
  x"6C",   x"90",   x"57",   x"AB",   x"1A",   x"E6",   x"21",   x"DD", 
  x"80",   x"7C",   x"BB",   x"47",   x"F6",   x"0A",   x"CD",   x"31", 
  x"77",   x"8B",   x"4C",   x"B0",   x"01",   x"FD",   x"3A",   x"C6", 
  x"9B",   x"67",   x"A0",   x"5C",   x"ED",   x"11",   x"D6",   x"2A", 
  x"5A",   x"A6",   x"61",   x"9D",   x"2C",   x"D0",   x"17",   x"EB", 
  x"B6",   x"4A",   x"8D",   x"71",   x"C0",   x"3C",   x"FB",   x"07", 
  x"41",   x"BD",   x"7A",   x"86",   x"37",   x"CB",   x"0C",   x"F0", 
  x"AD",   x"51",   x"96",   x"6A",   x"DB",   x"27",   x"E0",   x"1C", 
  x"D8",   x"24",   x"E3",   x"1F",   x"AE",   x"52",   x"95",   x"69", 
  x"34",   x"C8",   x"0F",   x"F3",   x"42",   x"BE",   x"79",   x"85", 
  x"C3",   x"3F",   x"F8",   x"04",   x"B5",   x"49",   x"8E",   x"72", 
  x"2F",   x"D3",   x"14",   x"E8",   x"59",   x"A5",   x"62",   x"9E", 
  x"EE",   x"12",   x"D5",   x"29",   x"98",   x"64",   x"A3",   x"5F", 
  x"02",   x"FE",   x"39",   x"C5",   x"74",   x"88",   x"4F",   x"B3", 
  x"F5",   x"09",   x"CE",   x"32",   x"83",   x"7F",   x"B8",   x"44", 
  x"19",   x"E5",   x"22",   x"DE",   x"6F",   x"93",   x"54",   x"A8", 
  x"B4",   x"48",   x"8F",   x"73",   x"C2",   x"3E",   x"F9",   x"05", 
  x"58",   x"A4",   x"63",   x"9F",   x"2E",   x"D2",   x"15",   x"E9", 
  x"AF",   x"53",   x"94",   x"68",   x"D9",   x"25",   x"E2",   x"1E", 
  x"43",   x"BF",   x"78",   x"84",   x"35",   x"C9",   x"0E",   x"F2", 
  x"82",   x"7E",   x"B9",   x"45",   x"F4",   x"08",   x"CF",   x"33", 
  x"6E",   x"92",   x"55",   x"A9",   x"18",   x"E4",   x"23",   x"DF", 
  x"99",   x"65",   x"A2",   x"5E",   x"EF",   x"13",   x"D4",   x"28", 
  x"75",   x"89",   x"4E",   x"B2",   x"03",   x"FF",   x"38",   x"C4", 
  x"00",   x"FD",   x"39",   x"C4",   x"72",   x"8F",   x"4B",   x"B6", 
  x"E4",   x"19",   x"DD",   x"20",   x"96",   x"6B",   x"AF",   x"52", 
  x"0B",   x"F6",   x"32",   x"CF",   x"79",   x"84",   x"40",   x"BD", 
  x"EF",   x"12",   x"D6",   x"2B",   x"9D",   x"60",   x"A4",   x"59", 
  x"16",   x"EB",   x"2F",   x"D2",   x"64",   x"99",   x"5D",   x"A0", 
  x"F2",   x"0F",   x"CB",   x"36",   x"80",   x"7D",   x"B9",   x"44", 
  x"1D",   x"E0",   x"24",   x"D9",   x"6F",   x"92",   x"56",   x"AB", 
  x"F9",   x"04",   x"C0",   x"3D",   x"8B",   x"76",   x"B2",   x"4F", 
  x"2C",   x"D1",   x"15",   x"E8",   x"5E",   x"A3",   x"67",   x"9A", 
  x"C8",   x"35",   x"F1",   x"0C",   x"BA",   x"47",   x"83",   x"7E", 
  x"27",   x"DA",   x"1E",   x"E3",   x"55",   x"A8",   x"6C",   x"91", 
  x"C3",   x"3E",   x"FA",   x"07",   x"B1",   x"4C",   x"88",   x"75", 
  x"3A",   x"C7",   x"03",   x"FE",   x"48",   x"B5",   x"71",   x"8C", 
  x"DE",   x"23",   x"E7",   x"1A",   x"AC",   x"51",   x"95",   x"68", 
  x"31",   x"CC",   x"08",   x"F5",   x"43",   x"BE",   x"7A",   x"87", 
  x"D5",   x"28",   x"EC",   x"11",   x"A7",   x"5A",   x"9E",   x"63", 
  x"58",   x"A5",   x"61",   x"9C",   x"2A",   x"D7",   x"13",   x"EE", 
  x"BC",   x"41",   x"85",   x"78",   x"CE",   x"33",   x"F7",   x"0A", 
  x"53",   x"AE",   x"6A",   x"97",   x"21",   x"DC",   x"18",   x"E5", 
  x"B7",   x"4A",   x"8E",   x"73",   x"C5",   x"38",   x"FC",   x"01", 
  x"4E",   x"B3",   x"77",   x"8A",   x"3C",   x"C1",   x"05",   x"F8", 
  x"AA",   x"57",   x"93",   x"6E",   x"D8",   x"25",   x"E1",   x"1C", 
  x"45",   x"B8",   x"7C",   x"81",   x"37",   x"CA",   x"0E",   x"F3", 
  x"A1",   x"5C",   x"98",   x"65",   x"D3",   x"2E",   x"EA",   x"17", 
  x"74",   x"89",   x"4D",   x"B0",   x"06",   x"FB",   x"3F",   x"C2", 
  x"90",   x"6D",   x"A9",   x"54",   x"E2",   x"1F",   x"DB",   x"26", 
  x"7F",   x"82",   x"46",   x"BB",   x"0D",   x"F0",   x"34",   x"C9", 
  x"9B",   x"66",   x"A2",   x"5F",   x"E9",   x"14",   x"D0",   x"2D", 
  x"62",   x"9F",   x"5B",   x"A6",   x"10",   x"ED",   x"29",   x"D4", 
  x"86",   x"7B",   x"BF",   x"42",   x"F4",   x"09",   x"CD",   x"30", 
  x"69",   x"94",   x"50",   x"AD",   x"1B",   x"E6",   x"22",   x"DF", 
  x"8D",   x"70",   x"B4",   x"49",   x"FF",   x"02",   x"C6",   x"3B", 
  x"00",   x"FE",   x"3F",   x"C1",   x"7E",   x"80",   x"41",   x"BF", 
  x"FC",   x"02",   x"C3",   x"3D",   x"82",   x"7C",   x"BD",   x"43", 
  x"3B",   x"C5",   x"04",   x"FA",   x"45",   x"BB",   x"7A",   x"84", 
  x"C7",   x"39",   x"F8",   x"06",   x"B9",   x"47",   x"86",   x"78", 
  x"76",   x"88",   x"49",   x"B7",   x"08",   x"F6",   x"37",   x"C9", 
  x"8A",   x"74",   x"B5",   x"4B",   x"F4",   x"0A",   x"CB",   x"35", 
  x"4D",   x"B3",   x"72",   x"8C",   x"33",   x"CD",   x"0C",   x"F2", 
  x"B1",   x"4F",   x"8E",   x"70",   x"CF",   x"31",   x"F0",   x"0E", 
  x"EC",   x"12",   x"D3",   x"2D",   x"92",   x"6C",   x"AD",   x"53", 
  x"10",   x"EE",   x"2F",   x"D1",   x"6E",   x"90",   x"51",   x"AF", 
  x"D7",   x"29",   x"E8",   x"16",   x"A9",   x"57",   x"96",   x"68", 
  x"2B",   x"D5",   x"14",   x"EA",   x"55",   x"AB",   x"6A",   x"94", 
  x"9A",   x"64",   x"A5",   x"5B",   x"E4",   x"1A",   x"DB",   x"25", 
  x"66",   x"98",   x"59",   x"A7",   x"18",   x"E6",   x"27",   x"D9", 
  x"A1",   x"5F",   x"9E",   x"60",   x"DF",   x"21",   x"E0",   x"1E", 
  x"5D",   x"A3",   x"62",   x"9C",   x"23",   x"DD",   x"1C",   x"E2", 
  x"1B",   x"E5",   x"24",   x"DA",   x"65",   x"9B",   x"5A",   x"A4", 
  x"E7",   x"19",   x"D8",   x"26",   x"99",   x"67",   x"A6",   x"58", 
  x"20",   x"DE",   x"1F",   x"E1",   x"5E",   x"A0",   x"61",   x"9F", 
  x"DC",   x"22",   x"E3",   x"1D",   x"A2",   x"5C",   x"9D",   x"63", 
  x"6D",   x"93",   x"52",   x"AC",   x"13",   x"ED",   x"2C",   x"D2", 
  x"91",   x"6F",   x"AE",   x"50",   x"EF",   x"11",   x"D0",   x"2E", 
  x"56",   x"A8",   x"69",   x"97",   x"28",   x"D6",   x"17",   x"E9", 
  x"AA",   x"54",   x"95",   x"6B",   x"D4",   x"2A",   x"EB",   x"15", 
  x"F7",   x"09",   x"C8",   x"36",   x"89",   x"77",   x"B6",   x"48", 
  x"0B",   x"F5",   x"34",   x"CA",   x"75",   x"8B",   x"4A",   x"B4", 
  x"CC",   x"32",   x"F3",   x"0D",   x"B2",   x"4C",   x"8D",   x"73", 
  x"30",   x"CE",   x"0F",   x"F1",   x"4E",   x"B0",   x"71",   x"8F", 
  x"81",   x"7F",   x"BE",   x"40",   x"FF",   x"01",   x"C0",   x"3E", 
  x"7D",   x"83",   x"42",   x"BC",   x"03",   x"FD",   x"3C",   x"C2", 
  x"BA",   x"44",   x"85",   x"7B",   x"C4",   x"3A",   x"FB",   x"05", 
  x"46",   x"B8",   x"79",   x"87",   x"38",   x"C6",   x"07",   x"F9", 
  x"00",   x"FF",   x"3D",   x"C2",   x"7A",   x"85",   x"47",   x"B8", 
  x"F4",   x"0B",   x"C9",   x"36",   x"8E",   x"71",   x"B3",   x"4C", 
  x"2B",   x"D4",   x"16",   x"E9",   x"51",   x"AE",   x"6C",   x"93", 
  x"DF",   x"20",   x"E2",   x"1D",   x"A5",   x"5A",   x"98",   x"67", 
  x"56",   x"A9",   x"6B",   x"94",   x"2C",   x"D3",   x"11",   x"EE", 
  x"A2",   x"5D",   x"9F",   x"60",   x"D8",   x"27",   x"E5",   x"1A", 
  x"7D",   x"82",   x"40",   x"BF",   x"07",   x"F8",   x"3A",   x"C5", 
  x"89",   x"76",   x"B4",   x"4B",   x"F3",   x"0C",   x"CE",   x"31", 
  x"AC",   x"53",   x"91",   x"6E",   x"D6",   x"29",   x"EB",   x"14", 
  x"58",   x"A7",   x"65",   x"9A",   x"22",   x"DD",   x"1F",   x"E0", 
  x"87",   x"78",   x"BA",   x"45",   x"FD",   x"02",   x"C0",   x"3F", 
  x"73",   x"8C",   x"4E",   x"B1",   x"09",   x"F6",   x"34",   x"CB", 
  x"FA",   x"05",   x"C7",   x"38",   x"80",   x"7F",   x"BD",   x"42", 
  x"0E",   x"F1",   x"33",   x"CC",   x"74",   x"8B",   x"49",   x"B6", 
  x"D1",   x"2E",   x"EC",   x"13",   x"AB",   x"54",   x"96",   x"69", 
  x"25",   x"DA",   x"18",   x"E7",   x"5F",   x"A0",   x"62",   x"9D", 
  x"9B",   x"64",   x"A6",   x"59",   x"E1",   x"1E",   x"DC",   x"23", 
  x"6F",   x"90",   x"52",   x"AD",   x"15",   x"EA",   x"28",   x"D7", 
  x"B0",   x"4F",   x"8D",   x"72",   x"CA",   x"35",   x"F7",   x"08", 
  x"44",   x"BB",   x"79",   x"86",   x"3E",   x"C1",   x"03",   x"FC", 
  x"CD",   x"32",   x"F0",   x"0F",   x"B7",   x"48",   x"8A",   x"75", 
  x"39",   x"C6",   x"04",   x"FB",   x"43",   x"BC",   x"7E",   x"81", 
  x"E6",   x"19",   x"DB",   x"24",   x"9C",   x"63",   x"A1",   x"5E", 
  x"12",   x"ED",   x"2F",   x"D0",   x"68",   x"97",   x"55",   x"AA", 
  x"37",   x"C8",   x"0A",   x"F5",   x"4D",   x"B2",   x"70",   x"8F", 
  x"C3",   x"3C",   x"FE",   x"01",   x"B9",   x"46",   x"84",   x"7B", 
  x"1C",   x"E3",   x"21",   x"DE",   x"66",   x"99",   x"5B",   x"A4", 
  x"E8",   x"17",   x"D5",   x"2A",   x"92",   x"6D",   x"AF",   x"50", 
  x"61",   x"9E",   x"5C",   x"A3",   x"1B",   x"E4",   x"26",   x"D9", 
  x"95",   x"6A",   x"A8",   x"57",   x"EF",   x"10",   x"D2",   x"2D", 
  x"4A",   x"B5",   x"77",   x"88",   x"30",   x"CF",   x"0D",   x"F2", 
  x"BE",   x"41",   x"83",   x"7C",   x"C4",   x"3B",   x"F9",   x"06" 
  );
  
end table_h_package;